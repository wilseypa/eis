--
--  Copyright (c) 2003 Launchbird Design Systems, Inc.
--  All rights reserved.
--  
--  Redistribution and use in source and binary forms, with or without modification, are permitted provided that the following conditions are met:
--    Redistributions of source code must retain the above copyright notice, this list of conditions and the following disclaimer.
--    Redistributions in binary form must reproduce the above copyright notice, this list of conditions and the following disclaimer in the documentation and/or other materials provided with the distribution.
--  
--  THIS SOFTWARE IS PROVIDED BY THE COPYRIGHT HOLDERS AND CONTRIBUTORS "AS IS" AND ANY EXPRESS OR IMPLIED WARRANTIES,
--  INCLUDING, BUT NOT LIMITED TO, THE IMPLIED WARRANTIES OF MERCHANTABILITY AND FITNESS FOR A PARTICULAR PURPOSE ARE DISCLAIMED.
--  IN NO EVENT SHALL THE COPYRIGHT OWNER OR CONTRIBUTORS BE LIABLE FOR ANY DIRECT, INDIRECT, INCIDENTAL, SPECIAL, EXEMPLARY,
--  OR CONSEQUENTIAL DAMAGES (INCLUDING, BUT NOT LIMITED TO, PROCUREMENT OF SUBSTITUTE GOODS OR SERVICES; LOSS OF USE, DATA, OR PROFITS;
--  OR BUSINESS INTERRUPTION) HOWEVER CAUSED AND ON ANY THEORY OF LIABILITY, WHETHER IN CONTRACT, STRICT LIABILITY, OR TORT
--  (INCLUDING NEGLIGENCE OR OTHERWISE) ARISING IN ANY WAY OUT OF THE USE OF THIS SOFTWARE, EVEN IF ADVISED OF THE POSSIBILITY OF SUCH DAMAGE.
--  
--  
--  Overview:
--  
--    Performs a radix 2 Fast Fourier Transform.
--    The FFT architecture is pipelined on a rank basis; each rank has its own butterfly and ranks are
--    isolated from each other using memory interleavers.  This FFT can perform calcualations on continuous
--    streaming data (one data set right after another).  More over, inputs and outputs are passed in pairs,
--    doubling the bandwidth.  For instance, a 2048 point FFT can perform a transform every 1024 cycles.
--  
--  Interface:
--  
--    Synchronization:
--      clock_c  : Clock input.
--      enable_i : Synchronous enable.
--      reset_i  : Synchronous reset.
--  
--    Inputs:
--      sync_i     : Input sync pulse must occur one frame prior to data input.
--      data_0_i   : Input data 0.  Width is 2 * precision.  Real on the left, imag on the right.
--      data_1_i   : Input data 1.  Width is 2 * precision.  Real on the left, imag on the right.
--  
--    Outputs:
--      sync_o     : Output sync pulse occurs one frame before data output.
--      data_0_o   : Output data 0.  Width is 2 * precision.  Real on the left, imag on the right.
--      data_1_o   : Output data 1.  Width is 2 * precision.  Real on the left, imag on the right.
--  
--  Built In Parameters:
--  
--    FFT Points   = 4096
--    Precision    = 18
--  
--  
--  
--  
--  Generated by Confluence 0.6.3  --  Launchbird Design Systems, Inc.  --  www.launchbird.com
--  
--  Build Date : Fri Aug 22 08:51:05 CDT 2003
--  
--  Interface
--  
--    Build Name    : cf_fft_4096_18
--    Clock Domains : clock_c  
--    Vector Input  : enable_i(1)
--    Vector Input  : reset_i(1)
--    Vector Input  : sync_i(1)
--    Vector Input  : data_0_i(36)
--    Vector Input  : data_1_i(36)
--    Vector Output : sync_o(1)
--    Vector Output : data_0_o(36)
--    Vector Output : data_1_o(36)
--  
--  
--  

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
entity cf_fft_4096_18_43 is
port (
clock_c : in std_logic;
i1 : in  unsigned(35 downto 0);
i2 : in  unsigned(35 downto 0);
i3 : in  unsigned(2 downto 0);
i4 : in  unsigned(0 downto 0);
i5 : in  unsigned(0 downto 0);
o1 : out unsigned(35 downto 0);
o2 : out unsigned(35 downto 0));
end entity cf_fft_4096_18_43;
architecture rtl of cf_fft_4096_18_43 is
signal n1 : unsigned(35 downto 0) := "000000000000000000000000000000000000";
signal n2 : unsigned(17 downto 0);
signal n3 : unsigned(17 downto 0);
signal n4 : unsigned(35 downto 0) := "000000000000000000000000000000000000";
signal n5 : unsigned(17 downto 0);
signal n6 : unsigned(17 downto 0);
signal n7 : unsigned(17 downto 0) := "000000000000000000";
signal n8 : unsigned(17 downto 0) := "000000000000000000";
signal n9 : unsigned(17 downto 0) := "000000000000000000";
signal n10 : unsigned(17 downto 0) := "000000000000000000";
signal n11 : unsigned(35 downto 0) := "000000000000000000000000000000000000";
signal n12 : unsigned(17 downto 0);
signal n13 : unsigned(17 downto 0);
signal n14 : unsigned(35 downto 0);
signal n15 : unsigned(17 downto 0);
signal n16 : unsigned(17 downto 0) := "000000000000000000";
signal n17 : unsigned(35 downto 0);
signal n18 : unsigned(17 downto 0);
signal n19 : unsigned(17 downto 0) := "000000000000000000";
signal n20 : unsigned(17 downto 0);
signal n21 : unsigned(17 downto 0) := "000000000000000000";
signal n22 : unsigned(35 downto 0);
signal n23 : unsigned(17 downto 0);
signal n24 : unsigned(17 downto 0) := "000000000000000000";
signal n25 : unsigned(35 downto 0);
signal n26 : unsigned(17 downto 0);
signal n27 : unsigned(17 downto 0) := "000000000000000000";
signal n28 : unsigned(17 downto 0);
signal n29 : unsigned(17 downto 0) := "000000000000000000";
signal n30 : unsigned(17 downto 0);
signal n31 : unsigned(17 downto 0);
signal n32 : unsigned(35 downto 0);
signal n33 : unsigned(35 downto 0) := "000000000000000000000000000000000000";
signal n34 : unsigned(17 downto 0);
signal n35 : unsigned(17 downto 0);
signal n36 : unsigned(35 downto 0);
signal n37 : unsigned(35 downto 0) := "000000000000000000000000000000000000";
begin
process (clock_c) begin
  if rising_edge(clock_c) then
    if i5 = "1" then
      n1 <= "000000000000000000000000000000000000";
    elsif i4 = "1" then
      n1 <= i1;
    end if;
  end if;
end process;
n2 <= n1(35 downto 35) &
  n1(34 downto 34) &
  n1(33 downto 33) &
  n1(32 downto 32) &
  n1(31 downto 31) &
  n1(30 downto 30) &
  n1(29 downto 29) &
  n1(28 downto 28) &
  n1(27 downto 27) &
  n1(26 downto 26) &
  n1(25 downto 25) &
  n1(24 downto 24) &
  n1(23 downto 23) &
  n1(22 downto 22) &
  n1(21 downto 21) &
  n1(20 downto 20) &
  n1(19 downto 19) &
  n1(18 downto 18);
n3 <= n1(17 downto 17) &
  n1(16 downto 16) &
  n1(15 downto 15) &
  n1(14 downto 14) &
  n1(13 downto 13) &
  n1(12 downto 12) &
  n1(11 downto 11) &
  n1(10 downto 10) &
  n1(9 downto 9) &
  n1(8 downto 8) &
  n1(7 downto 7) &
  n1(6 downto 6) &
  n1(5 downto 5) &
  n1(4 downto 4) &
  n1(3 downto 3) &
  n1(2 downto 2) &
  n1(1 downto 1) &
  n1(0 downto 0);
process (clock_c) begin
  if rising_edge(clock_c) then
    if i5 = "1" then
      n4 <= "000000000000000000000000000000000000";
    elsif i4 = "1" then
      n4 <= i2;
    end if;
  end if;
end process;
n5 <= n4(35 downto 35) &
  n4(34 downto 34) &
  n4(33 downto 33) &
  n4(32 downto 32) &
  n4(31 downto 31) &
  n4(30 downto 30) &
  n4(29 downto 29) &
  n4(28 downto 28) &
  n4(27 downto 27) &
  n4(26 downto 26) &
  n4(25 downto 25) &
  n4(24 downto 24) &
  n4(23 downto 23) &
  n4(22 downto 22) &
  n4(21 downto 21) &
  n4(20 downto 20) &
  n4(19 downto 19) &
  n4(18 downto 18);
n6 <= n4(17 downto 17) &
  n4(16 downto 16) &
  n4(15 downto 15) &
  n4(14 downto 14) &
  n4(13 downto 13) &
  n4(12 downto 12) &
  n4(11 downto 11) &
  n4(10 downto 10) &
  n4(9 downto 9) &
  n4(8 downto 8) &
  n4(7 downto 7) &
  n4(6 downto 6) &
  n4(5 downto 5) &
  n4(4 downto 4) &
  n4(3 downto 3) &
  n4(2 downto 2) &
  n4(1 downto 1) &
  n4(0 downto 0);
process (clock_c) begin
  if rising_edge(clock_c) then
    if i5 = "1" then
      n7 <= "000000000000000000";
    elsif i4 = "1" then
      n7 <= n2;
    end if;
  end if;
end process;
process (clock_c) begin
  if rising_edge(clock_c) then
    if i5 = "1" then
      n8 <= "000000000000000000";
    elsif i4 = "1" then
      n8 <= n7;
    end if;
  end if;
end process;
process (clock_c) begin
  if rising_edge(clock_c) then
    if i5 = "1" then
      n9 <= "000000000000000000";
    elsif i4 = "1" then
      n9 <= n3;
    end if;
  end if;
end process;
process (clock_c) begin
  if rising_edge(clock_c) then
    if i5 = "1" then
      n10 <= "000000000000000000";
    elsif i4 = "1" then
      n10 <= n9;
    end if;
  end if;
end process;
process (clock_c) begin
  if rising_edge(clock_c) then 
    if i4 = "1" then
      case i3 is
        when "000" => n11 <= "011111111111111111000000000000000000";
        when "001" => n11 <= "011101100100000110110011110000010000";
        when "010" => n11 <= "010110101000001001101001010111110110";
        when "011" => n11 <= "001100001111101111100010011011111001";
        when "100" => n11 <= "000000000000000000100000000000000000";
        when "101" => n11 <= "110011110000010000100010011011111001";
        when "110" => n11 <= "101001010111110110101001010111110110";
        when "111" => n11 <= "100010011011111001110011110000010000";
        when others => n11 <= "XXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX";
      end case;
    end if;
  end if;
end process;
n12 <= n11(35 downto 35) &
  n11(34 downto 34) &
  n11(33 downto 33) &
  n11(32 downto 32) &
  n11(31 downto 31) &
  n11(30 downto 30) &
  n11(29 downto 29) &
  n11(28 downto 28) &
  n11(27 downto 27) &
  n11(26 downto 26) &
  n11(25 downto 25) &
  n11(24 downto 24) &
  n11(23 downto 23) &
  n11(22 downto 22) &
  n11(21 downto 21) &
  n11(20 downto 20) &
  n11(19 downto 19) &
  n11(18 downto 18);
n13 <= n11(17 downto 17) &
  n11(16 downto 16) &
  n11(15 downto 15) &
  n11(14 downto 14) &
  n11(13 downto 13) &
  n11(12 downto 12) &
  n11(11 downto 11) &
  n11(10 downto 10) &
  n11(9 downto 9) &
  n11(8 downto 8) &
  n11(7 downto 7) &
  n11(6 downto 6) &
  n11(5 downto 5) &
  n11(4 downto 4) &
  n11(3 downto 3) &
  n11(2 downto 2) &
  n11(1 downto 1) &
  n11(0 downto 0);
n14 <= unsigned(signed(n5) * signed(n12));
n15 <= n14(34 downto 34) &
  n14(33 downto 33) &
  n14(32 downto 32) &
  n14(31 downto 31) &
  n14(30 downto 30) &
  n14(29 downto 29) &
  n14(28 downto 28) &
  n14(27 downto 27) &
  n14(26 downto 26) &
  n14(25 downto 25) &
  n14(24 downto 24) &
  n14(23 downto 23) &
  n14(22 downto 22) &
  n14(21 downto 21) &
  n14(20 downto 20) &
  n14(19 downto 19) &
  n14(18 downto 18) &
  n14(17 downto 17);
process (clock_c) begin
  if rising_edge(clock_c) then
    if i5 = "1" then
      n16 <= "000000000000000000";
    elsif i4 = "1" then
      n16 <= n15;
    end if;
  end if;
end process;
n17 <= unsigned(signed(n6) * signed(n13));
n18 <= n17(34 downto 34) &
  n17(33 downto 33) &
  n17(32 downto 32) &
  n17(31 downto 31) &
  n17(30 downto 30) &
  n17(29 downto 29) &
  n17(28 downto 28) &
  n17(27 downto 27) &
  n17(26 downto 26) &
  n17(25 downto 25) &
  n17(24 downto 24) &
  n17(23 downto 23) &
  n17(22 downto 22) &
  n17(21 downto 21) &
  n17(20 downto 20) &
  n17(19 downto 19) &
  n17(18 downto 18) &
  n17(17 downto 17);
process (clock_c) begin
  if rising_edge(clock_c) then
    if i5 = "1" then
      n19 <= "000000000000000000";
    elsif i4 = "1" then
      n19 <= n18;
    end if;
  end if;
end process;
n20 <= n16 - n19;
process (clock_c) begin
  if rising_edge(clock_c) then
    if i5 = "1" then
      n21 <= "000000000000000000";
    elsif i4 = "1" then
      n21 <= n20;
    end if;
  end if;
end process;
n22 <= unsigned(signed(n5) * signed(n13));
n23 <= n22(34 downto 34) &
  n22(33 downto 33) &
  n22(32 downto 32) &
  n22(31 downto 31) &
  n22(30 downto 30) &
  n22(29 downto 29) &
  n22(28 downto 28) &
  n22(27 downto 27) &
  n22(26 downto 26) &
  n22(25 downto 25) &
  n22(24 downto 24) &
  n22(23 downto 23) &
  n22(22 downto 22) &
  n22(21 downto 21) &
  n22(20 downto 20) &
  n22(19 downto 19) &
  n22(18 downto 18) &
  n22(17 downto 17);
process (clock_c) begin
  if rising_edge(clock_c) then
    if i5 = "1" then
      n24 <= "000000000000000000";
    elsif i4 = "1" then
      n24 <= n23;
    end if;
  end if;
end process;
n25 <= unsigned(signed(n6) * signed(n12));
n26 <= n25(34 downto 34) &
  n25(33 downto 33) &
  n25(32 downto 32) &
  n25(31 downto 31) &
  n25(30 downto 30) &
  n25(29 downto 29) &
  n25(28 downto 28) &
  n25(27 downto 27) &
  n25(26 downto 26) &
  n25(25 downto 25) &
  n25(24 downto 24) &
  n25(23 downto 23) &
  n25(22 downto 22) &
  n25(21 downto 21) &
  n25(20 downto 20) &
  n25(19 downto 19) &
  n25(18 downto 18) &
  n25(17 downto 17);
process (clock_c) begin
  if rising_edge(clock_c) then
    if i5 = "1" then
      n27 <= "000000000000000000";
    elsif i4 = "1" then
      n27 <= n26;
    end if;
  end if;
end process;
n28 <= n24 + n27;
process (clock_c) begin
  if rising_edge(clock_c) then
    if i5 = "1" then
      n29 <= "000000000000000000";
    elsif i4 = "1" then
      n29 <= n28;
    end if;
  end if;
end process;
n30 <= n8 + n21;
n31 <= n10 + n29;
n32 <= n30 & n31;
process (clock_c) begin
  if rising_edge(clock_c) then
    if i5 = "1" then
      n33 <= "000000000000000000000000000000000000";
    elsif i4 = "1" then
      n33 <= n32;
    end if;
  end if;
end process;
n34 <= n8 - n21;
n35 <= n10 - n29;
n36 <= n34 & n35;
process (clock_c) begin
  if rising_edge(clock_c) then
    if i5 = "1" then
      n37 <= "000000000000000000000000000000000000";
    elsif i4 = "1" then
      n37 <= n36;
    end if;
  end if;
end process;
o2 <= n37;
o1 <= n33;
end architecture rtl;

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
entity cf_fft_4096_18_42 is
port (
i1 : in  unsigned(0 downto 0);
i2 : in  unsigned(0 downto 0);
i3 : in  unsigned(0 downto 0);
i4 : in  unsigned(0 downto 0);
i5 : in  unsigned(2 downto 0);
o1 : out unsigned(0 downto 0));
end entity cf_fft_4096_18_42;
architecture rtl of cf_fft_4096_18_42 is
signal n1 : unsigned(2 downto 0);
signal n2 : unsigned(2 downto 0);
signal n3 : unsigned(2 downto 0);
signal n4 : unsigned(0 downto 0);
signal n5 : unsigned(0 downto 0);
signal n6 : unsigned(0 downto 0);
signal n7 : unsigned(0 downto 0);
signal n8 : unsigned(0 downto 0);
signal n9 : unsigned(0 downto 0);
begin
n1 <= "001";
n2 <= "011";
n3 <= "101";
n4 <= "1" when i5 = n1 else "0";
n5 <= "1" when i5 = n2 else "0";
n6 <= "1" when i5 = n3 else "0";
n7 <= i2 when n6 = "1" else i1;
n8 <= i3 when n5 = "1" else n7;
n9 <= i4 when n4 = "1" else n8;
o1 <= n9;
end architecture rtl;

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
entity cf_fft_4096_18_41 is
port (
i1 : in  unsigned(0 downto 0);
i2 : in  unsigned(0 downto 0);
i3 : in  unsigned(0 downto 0);
i4 : in  unsigned(0 downto 0);
i5 : in  unsigned(0 downto 0);
i6 : in  unsigned(0 downto 0);
i7 : in  unsigned(0 downto 0);
i8 : in  unsigned(2 downto 0);
o1 : out unsigned(0 downto 0));
end entity cf_fft_4096_18_41;
architecture rtl of cf_fft_4096_18_41 is
signal n1 : unsigned(2 downto 0);
signal n2 : unsigned(2 downto 0);
signal n3 : unsigned(2 downto 0);
signal n4 : unsigned(0 downto 0);
signal n5 : unsigned(0 downto 0);
signal n6 : unsigned(0 downto 0);
signal n7 : unsigned(0 downto 0);
signal n8 : unsigned(0 downto 0);
signal n9 : unsigned(0 downto 0);
signal s10_1 : unsigned(0 downto 0);
component cf_fft_4096_18_42 is
port (
i1 : in  unsigned(0 downto 0);
i2 : in  unsigned(0 downto 0);
i3 : in  unsigned(0 downto 0);
i4 : in  unsigned(0 downto 0);
i5 : in  unsigned(2 downto 0);
o1 : out unsigned(0 downto 0));
end component cf_fft_4096_18_42;
begin
n1 <= "010";
n2 <= "100";
n3 <= "110";
n4 <= "1" when i8 = n1 else "0";
n5 <= "1" when i8 = n2 else "0";
n6 <= "1" when i8 = n3 else "0";
n7 <= i5 when n6 = "1" else s10_1;
n8 <= i6 when n5 = "1" else n7;
n9 <= i7 when n4 = "1" else n8;
s10 : cf_fft_4096_18_42 port map (i1, i2, i3, i4, i8, s10_1);
o1 <= n9;
end architecture rtl;

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
entity cf_fft_4096_18_40 is
port (
o1 : out unsigned(0 downto 0);
o2 : out unsigned(0 downto 0);
o3 : out unsigned(0 downto 0);
o4 : out unsigned(0 downto 0);
o5 : out unsigned(0 downto 0);
o6 : out unsigned(0 downto 0);
o7 : out unsigned(0 downto 0);
o8 : out unsigned(0 downto 0));
end entity cf_fft_4096_18_40;
architecture rtl of cf_fft_4096_18_40 is
signal n1 : unsigned(0 downto 0);
signal n2 : unsigned(0 downto 0);
signal n3 : unsigned(0 downto 0);
signal n4 : unsigned(0 downto 0);
signal n5 : unsigned(0 downto 0);
signal n6 : unsigned(0 downto 0);
signal n7 : unsigned(0 downto 0);
signal n8 : unsigned(0 downto 0);
begin
n1 <= "0";
n2 <= "1";
n3 <= "0";
n4 <= "1";
n5 <= "0";
n6 <= "1";
n7 <= "0";
n8 <= "0";
o8 <= n8;
o7 <= n7;
o6 <= n6;
o5 <= n5;
o4 <= n4;
o3 <= n3;
o2 <= n2;
o1 <= n1;
end architecture rtl;

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
entity cf_fft_4096_18_39 is
port (
i1 : in  unsigned(0 downto 0);
i2 : in  unsigned(0 downto 0);
i3 : in  unsigned(0 downto 0);
i4 : in  unsigned(2 downto 0);
o1 : out unsigned(0 downto 0));
end entity cf_fft_4096_18_39;
architecture rtl of cf_fft_4096_18_39 is
signal n1 : unsigned(2 downto 0);
signal n2 : unsigned(2 downto 0);
signal n3 : unsigned(2 downto 0);
signal n4 : unsigned(0 downto 0);
signal n5 : unsigned(0 downto 0);
signal n6 : unsigned(0 downto 0);
signal n7 : unsigned(0 downto 0);
signal n8 : unsigned(0 downto 0);
signal n9 : unsigned(0 downto 0);
signal n10 : unsigned(0 downto 0);
begin
n1 <= "010";
n2 <= "100";
n3 <= "110";
n4 <= "1" when i4 = n1 else "0";
n5 <= "1" when i4 = n2 else "0";
n6 <= "1" when i4 = n3 else "0";
n7 <= i1 when n6 = "1" else n10;
n8 <= i2 when n5 = "1" else n7;
n9 <= i3 when n4 = "1" else n8;
n10 <= "1";
o1 <= n9;
end architecture rtl;

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
entity cf_fft_4096_18_38 is
port (
i1 : in  unsigned(2 downto 0);
o1 : out unsigned(0 downto 0));
end entity cf_fft_4096_18_38;
architecture rtl of cf_fft_4096_18_38 is
signal n1 : unsigned(0 downto 0);
signal n2 : unsigned(0 downto 0);
signal n3 : unsigned(0 downto 0);
signal n4 : unsigned(0 downto 0);
signal n5 : unsigned(2 downto 0);
signal n6 : unsigned(0 downto 0);
signal n7 : unsigned(0 downto 0);
signal s8_1 : unsigned(0 downto 0);
component cf_fft_4096_18_39 is
port (
i1 : in  unsigned(0 downto 0);
i2 : in  unsigned(0 downto 0);
i3 : in  unsigned(0 downto 0);
i4 : in  unsigned(2 downto 0);
o1 : out unsigned(0 downto 0));
end component cf_fft_4096_18_39;
begin
n1 <= "0";
n2 <= "0";
n3 <= "0";
n4 <= "0";
n5 <= "000";
n6 <= "1" when i1 = n5 else "0";
n7 <= n4 when n6 = "1" else s8_1;
s8 : cf_fft_4096_18_39 port map (n1, n2, n3, i1, s8_1);
o1 <= n7;
end architecture rtl;

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
entity cf_fft_4096_18_37 is
port (
clock_c : in std_logic;
i1 : in  unsigned(1 downto 0);
i2 : in  unsigned(0 downto 0);
i3 : in  unsigned(0 downto 0);
o1 : out unsigned(0 downto 0));
end entity cf_fft_4096_18_37;
architecture rtl of cf_fft_4096_18_37 is
signal n1 : unsigned(2 downto 0);
signal n2 : unsigned(2 downto 0);
signal n3 : unsigned(0 downto 0);
signal n4 : unsigned(0 downto 0);
signal n5 : unsigned(0 downto 0) := "0";
signal s6_1 : unsigned(0 downto 0);
signal s7_1 : unsigned(0 downto 0);
signal s7_2 : unsigned(0 downto 0);
signal s7_3 : unsigned(0 downto 0);
signal s7_4 : unsigned(0 downto 0);
signal s7_5 : unsigned(0 downto 0);
signal s7_6 : unsigned(0 downto 0);
signal s7_7 : unsigned(0 downto 0);
signal s7_8 : unsigned(0 downto 0);
signal s8_1 : unsigned(0 downto 0);
component cf_fft_4096_18_41 is
port (
i1 : in  unsigned(0 downto 0);
i2 : in  unsigned(0 downto 0);
i3 : in  unsigned(0 downto 0);
i4 : in  unsigned(0 downto 0);
i5 : in  unsigned(0 downto 0);
i6 : in  unsigned(0 downto 0);
i7 : in  unsigned(0 downto 0);
i8 : in  unsigned(2 downto 0);
o1 : out unsigned(0 downto 0));
end component cf_fft_4096_18_41;
component cf_fft_4096_18_40 is
port (
o1 : out unsigned(0 downto 0);
o2 : out unsigned(0 downto 0);
o3 : out unsigned(0 downto 0);
o4 : out unsigned(0 downto 0);
o5 : out unsigned(0 downto 0);
o6 : out unsigned(0 downto 0);
o7 : out unsigned(0 downto 0);
o8 : out unsigned(0 downto 0));
end component cf_fft_4096_18_40;
component cf_fft_4096_18_38 is
port (
i1 : in  unsigned(2 downto 0);
o1 : out unsigned(0 downto 0));
end component cf_fft_4096_18_38;
begin
n1 <= "000";
n2 <= i1 & n5;
n3 <= "1" when n2 = n1 else "0";
n4 <= s7_8 when n3 = "1" else s6_1;
process (clock_c) begin
  if rising_edge(clock_c) then
    if i3 = "1" then
      n5 <= "0";
    elsif i2 = "1" then
      n5 <= n4;
    end if;
  end if;
end process;
s6 : cf_fft_4096_18_41 port map (s7_1, s7_2, s7_3, s7_4, s7_5, s7_6, s7_7, n2, s6_1);
s7 : cf_fft_4096_18_40 port map (s7_1, s7_2, s7_3, s7_4, s7_5, s7_6, s7_7, s7_8);
s8 : cf_fft_4096_18_38 port map (n2, s8_1);
o1 <= s8_1;
end architecture rtl;

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
entity cf_fft_4096_18_36 is
port (
i1 : in  unsigned(0 downto 0);
i2 : in  unsigned(0 downto 0);
i3 : in  unsigned(0 downto 0);
i4 : in  unsigned(0 downto 0);
i5 : in  unsigned(1 downto 0);
o1 : out unsigned(0 downto 0));
end entity cf_fft_4096_18_36;
architecture rtl of cf_fft_4096_18_36 is
signal n1 : unsigned(1 downto 0);
signal n2 : unsigned(1 downto 0);
signal n3 : unsigned(1 downto 0);
signal n4 : unsigned(0 downto 0);
signal n5 : unsigned(0 downto 0);
signal n6 : unsigned(0 downto 0);
signal n7 : unsigned(0 downto 0);
signal n8 : unsigned(0 downto 0);
signal n9 : unsigned(0 downto 0);
begin
n1 <= "00";
n2 <= "10";
n3 <= "01";
n4 <= "1" when i5 = n1 else "0";
n5 <= "1" when i5 = n2 else "0";
n6 <= "1" when i5 = n3 else "0";
n7 <= i2 when n6 = "1" else i1;
n8 <= i3 when n5 = "1" else n7;
n9 <= i4 when n4 = "1" else n8;
o1 <= n9;
end architecture rtl;

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
entity cf_fft_4096_18_35 is
port (
i1 : in  unsigned(1 downto 0);
o1 : out unsigned(0 downto 0));
end entity cf_fft_4096_18_35;
architecture rtl of cf_fft_4096_18_35 is
signal n1 : unsigned(0 downto 0);
signal n2 : unsigned(0 downto 0);
signal n3 : unsigned(1 downto 0);
signal n4 : unsigned(1 downto 0);
signal n5 : unsigned(0 downto 0);
signal n6 : unsigned(0 downto 0);
signal n7 : unsigned(0 downto 0);
signal n8 : unsigned(0 downto 0);
signal n9 : unsigned(0 downto 0);
begin
n1 <= "0";
n2 <= "0";
n3 <= "00";
n4 <= "10";
n5 <= "1" when i1 = n3 else "0";
n6 <= "1" when i1 = n4 else "0";
n7 <= n1 when n6 = "1" else n9;
n8 <= n2 when n5 = "1" else n7;
n9 <= "1";
o1 <= n8;
end architecture rtl;

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
entity cf_fft_4096_18_34 is
port (
clock_c : in std_logic;
i1 : in  unsigned(0 downto 0);
i2 : in  unsigned(0 downto 0);
i3 : in  unsigned(0 downto 0);
o1 : out unsigned(0 downto 0));
end entity cf_fft_4096_18_34;
architecture rtl of cf_fft_4096_18_34 is
signal n1 : unsigned(0 downto 0);
signal n2 : unsigned(0 downto 0);
signal n3 : unsigned(0 downto 0);
signal n4 : unsigned(0 downto 0);
signal n5 : unsigned(1 downto 0);
signal n6 : unsigned(0 downto 0) := "0";
signal s7_1 : unsigned(0 downto 0);
signal s8_1 : unsigned(0 downto 0);
component cf_fft_4096_18_36 is
port (
i1 : in  unsigned(0 downto 0);
i2 : in  unsigned(0 downto 0);
i3 : in  unsigned(0 downto 0);
i4 : in  unsigned(0 downto 0);
i5 : in  unsigned(1 downto 0);
o1 : out unsigned(0 downto 0));
end component cf_fft_4096_18_36;
component cf_fft_4096_18_35 is
port (
i1 : in  unsigned(1 downto 0);
o1 : out unsigned(0 downto 0));
end component cf_fft_4096_18_35;
begin
n1 <= "0";
n2 <= "1";
n3 <= "1";
n4 <= "0";
n5 <= i1 & n6;
process (clock_c) begin
  if rising_edge(clock_c) then
    if i3 = "1" then
      n6 <= "0";
    elsif i2 = "1" then
      n6 <= s7_1;
    end if;
  end if;
end process;
s7 : cf_fft_4096_18_36 port map (n1, n2, n3, n4, n5, s7_1);
s8 : cf_fft_4096_18_35 port map (n5, s8_1);
o1 <= s8_1;
end architecture rtl;

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
entity cf_fft_4096_18_33 is
port (
clock_c : in std_logic;
i1 : in  unsigned(71 downto 0);
i2 : in  unsigned(0 downto 0);
i3 : in  unsigned(9 downto 0);
i4 : in  unsigned(0 downto 0);
i5 : in  unsigned(0 downto 0);
i6 : in  unsigned(0 downto 0);
o1 : out unsigned(71 downto 0));
end entity cf_fft_4096_18_33;
architecture rtl of cf_fft_4096_18_33 is
signal n1 : unsigned(9 downto 0);
signal n2 : unsigned(9 downto 0);
signal n3 : unsigned(9 downto 0) := "0000000000";
signal n4 : unsigned(0 downto 0);
signal n5 : unsigned(0 downto 0);
signal n6 : unsigned(71 downto 0);
signal n6a : unsigned(9 downto 0) := "0000000000";
type   n6mt is array (1023 downto 0) of unsigned(71 downto 0);
signal n6m : n6mt;
signal n7 : unsigned(0 downto 0);
signal n8 : unsigned(71 downto 0);
signal n8a : unsigned(9 downto 0) := "0000000000";
type   n8mt is array (1023 downto 0) of unsigned(71 downto 0);
signal n8m : n8mt;
signal n9 : unsigned(0 downto 0) := "0";
signal n10 : unsigned(71 downto 0);
signal n11 : unsigned(0 downto 0);
signal s12_1 : unsigned(0 downto 0);
component cf_fft_4096_18_34 is
port (
clock_c : in std_logic;
i1 : in  unsigned(0 downto 0);
i2 : in  unsigned(0 downto 0);
i3 : in  unsigned(0 downto 0);
o1 : out unsigned(0 downto 0));
end component cf_fft_4096_18_34;
begin
n1 <= "0000000001";
n2 <= n3 + n1;
process (clock_c) begin
  if rising_edge(clock_c) then
    if n11 = "1" then
      n3 <= "0000000000";
    elsif i5 = "1" then
      n3 <= n2;
    end if;
  end if;
end process;
n4 <= not s12_1;
n5 <= i4 and n4;
process (clock_c) begin
  if rising_edge(clock_c) then
    if i5 = "1" then
      if n5 = "1" then
        n6m(to_integer(i3)) <= i1;
      end if;
      n6a <= n3;
    end if;
  end if;
end process;
n6 <= n6m(to_integer(n6a));
n7 <= i4 and s12_1;
process (clock_c) begin
  if rising_edge(clock_c) then
    if i5 = "1" then
      if n7 = "1" then
        n8m(to_integer(i3)) <= i1;
      end if;
      n8a <= n3;
    end if;
  end if;
end process;
n8 <= n8m(to_integer(n8a));
process (clock_c) begin
  if rising_edge(clock_c) then
    if i6 = "1" then
      n9 <= "0";
    elsif i5 = "1" then
      n9 <= n4;
    end if;
  end if;
end process;
n10 <= n8 when n9 = "1" else n6;
n11 <= i2 or i6;
s12 : cf_fft_4096_18_34 port map (clock_c, i2, i5, i6, s12_1);
o1 <= n10;
end architecture rtl;

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
entity cf_fft_4096_18_32 is
port (
clock_c : in std_logic;
i1 : in  unsigned(71 downto 0);
i2 : in  unsigned(0 downto 0);
i3 : in  unsigned(9 downto 0);
i4 : in  unsigned(0 downto 0);
i5 : in  unsigned(0 downto 0);
i6 : in  unsigned(0 downto 0);
o1 : out unsigned(0 downto 0);
o2 : out unsigned(0 downto 0);
o3 : out unsigned(71 downto 0));
end entity cf_fft_4096_18_32;
architecture rtl of cf_fft_4096_18_32 is
signal n1 : unsigned(9 downto 0);
signal n2 : unsigned(9 downto 0);
signal n3 : unsigned(9 downto 0) := "0000000000";
signal n4 : unsigned(0 downto 0);
signal n5 : unsigned(0 downto 0) := "0";
signal n6 : unsigned(9 downto 0);
signal n7 : unsigned(0 downto 0);
signal n8 : unsigned(0 downto 0);
signal n9 : unsigned(71 downto 0);
signal n9a : unsigned(9 downto 0) := "0000000000";
type   n9mt is array (1023 downto 0) of unsigned(71 downto 0);
signal n9m : n9mt;
signal n10 : unsigned(0 downto 0);
signal n11 : unsigned(71 downto 0);
signal n11a : unsigned(9 downto 0) := "0000000000";
type   n11mt is array (1023 downto 0) of unsigned(71 downto 0);
signal n11m : n11mt;
signal n12 : unsigned(0 downto 0) := "0";
signal n13 : unsigned(71 downto 0);
signal n14 : unsigned(0 downto 0);
signal s15_1 : unsigned(0 downto 0);
component cf_fft_4096_18_34 is
port (
clock_c : in std_logic;
i1 : in  unsigned(0 downto 0);
i2 : in  unsigned(0 downto 0);
i3 : in  unsigned(0 downto 0);
o1 : out unsigned(0 downto 0));
end component cf_fft_4096_18_34;
begin
n1 <= "0000000001";
n2 <= n3 + n1;
process (clock_c) begin
  if rising_edge(clock_c) then
    if n14 = "1" then
      n3 <= "0000000000";
    elsif i5 = "1" then
      n3 <= n2;
    end if;
  end if;
end process;
n4 <= not s15_1;
process (clock_c) begin
  if rising_edge(clock_c) then
    if i6 = "1" then
      n5 <= "0";
    elsif i5 = "1" then
      n5 <= i2;
    end if;
  end if;
end process;
n6 <= "0000000000";
n7 <= "1" when n3 = n6 else "0";
n8 <= i4 and n4;
process (clock_c) begin
  if rising_edge(clock_c) then
    if i5 = "1" then
      if n8 = "1" then
        n9m(to_integer(i3)) <= i1;
      end if;
      n9a <= n3;
    end if;
  end if;
end process;
n9 <= n9m(to_integer(n9a));
n10 <= i4 and s15_1;
process (clock_c) begin
  if rising_edge(clock_c) then
    if i5 = "1" then
      if n10 = "1" then
        n11m(to_integer(i3)) <= i1;
      end if;
      n11a <= n3;
    end if;
  end if;
end process;
n11 <= n11m(to_integer(n11a));
process (clock_c) begin
  if rising_edge(clock_c) then
    if i6 = "1" then
      n12 <= "0";
    elsif i5 = "1" then
      n12 <= n4;
    end if;
  end if;
end process;
n13 <= n11 when n12 = "1" else n9;
n14 <= i2 or i6;
s15 : cf_fft_4096_18_34 port map (clock_c, i2, i5, i6, s15_1);
o3 <= n13;
o2 <= n7;
o1 <= n5;
end architecture rtl;

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
entity cf_fft_4096_18_31 is
port (
i1 : in  unsigned(0 downto 0);
i2 : in  unsigned(0 downto 0);
i3 : in  unsigned(0 downto 0);
i4 : in  unsigned(2 downto 0);
o1 : out unsigned(0 downto 0));
end entity cf_fft_4096_18_31;
architecture rtl of cf_fft_4096_18_31 is
signal n1 : unsigned(2 downto 0);
signal n2 : unsigned(2 downto 0);
signal n3 : unsigned(2 downto 0);
signal n4 : unsigned(0 downto 0);
signal n5 : unsigned(0 downto 0);
signal n6 : unsigned(0 downto 0);
signal n7 : unsigned(0 downto 0);
signal n8 : unsigned(0 downto 0);
signal n9 : unsigned(0 downto 0);
signal n10 : unsigned(0 downto 0);
begin
n1 <= "110";
n2 <= "001";
n3 <= "011";
n4 <= "1" when i4 = n1 else "0";
n5 <= "1" when i4 = n2 else "0";
n6 <= "1" when i4 = n3 else "0";
n7 <= i1 when n6 = "1" else n10;
n8 <= i2 when n5 = "1" else n7;
n9 <= i3 when n4 = "1" else n8;
n10 <= "1";
o1 <= n9;
end architecture rtl;

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
entity cf_fft_4096_18_30 is
port (
i1 : in  unsigned(0 downto 0);
i2 : in  unsigned(0 downto 0);
i3 : in  unsigned(0 downto 0);
i4 : in  unsigned(0 downto 0);
i5 : in  unsigned(0 downto 0);
i6 : in  unsigned(0 downto 0);
i7 : in  unsigned(2 downto 0);
o1 : out unsigned(0 downto 0));
end entity cf_fft_4096_18_30;
architecture rtl of cf_fft_4096_18_30 is
signal n1 : unsigned(2 downto 0);
signal n2 : unsigned(2 downto 0);
signal n3 : unsigned(2 downto 0);
signal n4 : unsigned(0 downto 0);
signal n5 : unsigned(0 downto 0);
signal n6 : unsigned(0 downto 0);
signal n7 : unsigned(0 downto 0);
signal n8 : unsigned(0 downto 0);
signal n9 : unsigned(0 downto 0);
signal s10_1 : unsigned(0 downto 0);
component cf_fft_4096_18_31 is
port (
i1 : in  unsigned(0 downto 0);
i2 : in  unsigned(0 downto 0);
i3 : in  unsigned(0 downto 0);
i4 : in  unsigned(2 downto 0);
o1 : out unsigned(0 downto 0));
end component cf_fft_4096_18_31;
begin
n1 <= "000";
n2 <= "010";
n3 <= "100";
n4 <= "1" when i7 = n1 else "0";
n5 <= "1" when i7 = n2 else "0";
n6 <= "1" when i7 = n3 else "0";
n7 <= i4 when n6 = "1" else s10_1;
n8 <= i5 when n5 = "1" else n7;
n9 <= i6 when n4 = "1" else n8;
s10 : cf_fft_4096_18_31 port map (i1, i2, i3, i7, s10_1);
o1 <= n9;
end architecture rtl;

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
entity cf_fft_4096_18_29 is
port (
clock_c : in std_logic;
i1 : in  unsigned(1 downto 0);
i2 : in  unsigned(0 downto 0);
i3 : in  unsigned(0 downto 0);
o1 : out unsigned(0 downto 0));
end entity cf_fft_4096_18_29;
architecture rtl of cf_fft_4096_18_29 is
signal n1 : unsigned(0 downto 0);
signal n2 : unsigned(0 downto 0);
signal n3 : unsigned(0 downto 0);
signal n4 : unsigned(0 downto 0);
signal n5 : unsigned(0 downto 0);
signal n6 : unsigned(0 downto 0);
signal n7 : unsigned(0 downto 0);
signal n8 : unsigned(0 downto 0);
signal n9 : unsigned(0 downto 0);
signal n10 : unsigned(0 downto 0);
signal n11 : unsigned(0 downto 0);
signal n12 : unsigned(0 downto 0);
signal n13 : unsigned(2 downto 0);
signal n14 : unsigned(0 downto 0) := "0";
signal s15_1 : unsigned(0 downto 0);
signal s16_1 : unsigned(0 downto 0);
component cf_fft_4096_18_30 is
port (
i1 : in  unsigned(0 downto 0);
i2 : in  unsigned(0 downto 0);
i3 : in  unsigned(0 downto 0);
i4 : in  unsigned(0 downto 0);
i5 : in  unsigned(0 downto 0);
i6 : in  unsigned(0 downto 0);
i7 : in  unsigned(2 downto 0);
o1 : out unsigned(0 downto 0));
end component cf_fft_4096_18_30;
begin
n1 <= "0";
n2 <= "1";
n3 <= "1";
n4 <= "1";
n5 <= "0";
n6 <= "0";
n7 <= "0";
n8 <= "1";
n9 <= "1";
n10 <= "1";
n11 <= "0";
n12 <= "0";
n13 <= i1 & n14;
process (clock_c) begin
  if rising_edge(clock_c) then
    if i3 = "1" then
      n14 <= "0";
    elsif i2 = "1" then
      n14 <= s15_1;
    end if;
  end if;
end process;
s15 : cf_fft_4096_18_30 port map (n1, n2, n3, n4, n5, n6, n13, s15_1);
s16 : cf_fft_4096_18_30 port map (n7, n8, n9, n10, n11, n12, n13, s16_1);
o1 <= s16_1;
end architecture rtl;

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
entity cf_fft_4096_18_28 is
port (
clock_c : in std_logic;
i1 : in  unsigned(0 downto 0);
i2 : in  unsigned(0 downto 0);
i3 : in  unsigned(0 downto 0);
o1 : out unsigned(10 downto 0);
o2 : out unsigned(0 downto 0));
end entity cf_fft_4096_18_28;
architecture rtl of cf_fft_4096_18_28 is
signal n1 : unsigned(10 downto 0);
signal n2 : unsigned(10 downto 0);
signal n3 : unsigned(10 downto 0) := "00000000000";
signal n4 : unsigned(10 downto 0);
signal n5 : unsigned(0 downto 0);
signal n6 : unsigned(1 downto 0);
signal n7 : unsigned(0 downto 0) := "0";
signal n8 : unsigned(0 downto 0);
signal n9 : unsigned(0 downto 0);
signal n10 : unsigned(0 downto 0);
signal s11_1 : unsigned(0 downto 0);
component cf_fft_4096_18_29 is
port (
clock_c : in std_logic;
i1 : in  unsigned(1 downto 0);
i2 : in  unsigned(0 downto 0);
i3 : in  unsigned(0 downto 0);
o1 : out unsigned(0 downto 0));
end component cf_fft_4096_18_29;
begin
n1 <= "00000000001";
n2 <= n3 + n1;
process (clock_c) begin
  if rising_edge(clock_c) then
    if n9 = "1" then
      n3 <= "00000000000";
    elsif n10 = "1" then
      n3 <= n2;
    end if;
  end if;
end process;
n4 <= "11111111111";
n5 <= "1" when n3 = n4 else "0";
n6 <= i1 & n5;
process (clock_c) begin
  if rising_edge(clock_c) then
    if i3 = "1" then
      n7 <= "0";
    elsif i2 = "1" then
      n7 <= s11_1;
    end if;
  end if;
end process;
n8 <= n7 and n5;
n9 <= i1 or i3;
n10 <= s11_1 and i2;
s11 : cf_fft_4096_18_29 port map (clock_c, n6, i2, i3, s11_1);
o2 <= n8;
o1 <= n3;
end architecture rtl;

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
entity cf_fft_4096_18_27 is
port (
clock_c : in std_logic;
i1 : in  unsigned(0 downto 0);
i2 : in  unsigned(35 downto 0);
i3 : in  unsigned(35 downto 0);
i4 : in  unsigned(0 downto 0);
i5 : in  unsigned(0 downto 0);
o1 : out unsigned(0 downto 0);
o2 : out unsigned(35 downto 0);
o3 : out unsigned(35 downto 0));
end entity cf_fft_4096_18_27;
architecture rtl of cf_fft_4096_18_27 is
signal n1 : unsigned(2 downto 0);
signal n2 : unsigned(71 downto 0);
signal n3 : unsigned(0 downto 0) := "0";
signal n4 : unsigned(0 downto 0) := "0";
signal n5 : unsigned(0 downto 0) := "0";
signal n6 : unsigned(0 downto 0) := "0";
signal n7 : unsigned(9 downto 0);
signal n8 : unsigned(9 downto 0) := "0000000000";
signal n9 : unsigned(9 downto 0) := "0000000000";
signal n10 : unsigned(9 downto 0) := "0000000000";
signal n11 : unsigned(9 downto 0) := "0000000000";
signal n12 : unsigned(0 downto 0);
signal n13 : unsigned(0 downto 0) := "0";
signal n14 : unsigned(0 downto 0) := "0";
signal n15 : unsigned(0 downto 0) := "0";
signal n16 : unsigned(0 downto 0) := "0";
signal n17 : unsigned(0 downto 0);
signal n18 : unsigned(1 downto 0);
signal n19 : unsigned(35 downto 0);
signal n20 : unsigned(35 downto 0);
signal n21 : unsigned(35 downto 0);
signal n22 : unsigned(35 downto 0);
signal n23 : unsigned(35 downto 0);
signal n24 : unsigned(35 downto 0);
signal s25_1 : unsigned(35 downto 0);
signal s25_2 : unsigned(35 downto 0);
signal s26_1 : unsigned(0 downto 0);
signal s27_1 : unsigned(71 downto 0);
signal s28_1 : unsigned(0 downto 0);
signal s28_2 : unsigned(0 downto 0);
signal s28_3 : unsigned(71 downto 0);
signal s29_1 : unsigned(10 downto 0);
signal s29_2 : unsigned(0 downto 0);
component cf_fft_4096_18_43 is
port (
clock_c : in std_logic;
i1 : in  unsigned(35 downto 0);
i2 : in  unsigned(35 downto 0);
i3 : in  unsigned(2 downto 0);
i4 : in  unsigned(0 downto 0);
i5 : in  unsigned(0 downto 0);
o1 : out unsigned(35 downto 0);
o2 : out unsigned(35 downto 0));
end component cf_fft_4096_18_43;
component cf_fft_4096_18_37 is
port (
clock_c : in std_logic;
i1 : in  unsigned(1 downto 0);
i2 : in  unsigned(0 downto 0);
i3 : in  unsigned(0 downto 0);
o1 : out unsigned(0 downto 0));
end component cf_fft_4096_18_37;
component cf_fft_4096_18_33 is
port (
clock_c : in std_logic;
i1 : in  unsigned(71 downto 0);
i2 : in  unsigned(0 downto 0);
i3 : in  unsigned(9 downto 0);
i4 : in  unsigned(0 downto 0);
i5 : in  unsigned(0 downto 0);
i6 : in  unsigned(0 downto 0);
o1 : out unsigned(71 downto 0));
end component cf_fft_4096_18_33;
component cf_fft_4096_18_32 is
port (
clock_c : in std_logic;
i1 : in  unsigned(71 downto 0);
i2 : in  unsigned(0 downto 0);
i3 : in  unsigned(9 downto 0);
i4 : in  unsigned(0 downto 0);
i5 : in  unsigned(0 downto 0);
i6 : in  unsigned(0 downto 0);
o1 : out unsigned(0 downto 0);
o2 : out unsigned(0 downto 0);
o3 : out unsigned(71 downto 0));
end component cf_fft_4096_18_32;
component cf_fft_4096_18_28 is
port (
clock_c : in std_logic;
i1 : in  unsigned(0 downto 0);
i2 : in  unsigned(0 downto 0);
i3 : in  unsigned(0 downto 0);
o1 : out unsigned(10 downto 0);
o2 : out unsigned(0 downto 0));
end component cf_fft_4096_18_28;
begin
n1 <= s29_1(10 downto 10) &
  s29_1(9 downto 9) &
  s29_1(8 downto 8);
n2 <= s25_1 & s25_2;
process (clock_c) begin
  if rising_edge(clock_c) then
    if i5 = "1" then
      n3 <= "0";
    elsif i4 = "1" then
      n3 <= s29_2;
    end if;
  end if;
end process;
process (clock_c) begin
  if rising_edge(clock_c) then
    if i5 = "1" then
      n4 <= "0";
    elsif i4 = "1" then
      n4 <= n3;
    end if;
  end if;
end process;
process (clock_c) begin
  if rising_edge(clock_c) then
    if i5 = "1" then
      n5 <= "0";
    elsif i4 = "1" then
      n5 <= n4;
    end if;
  end if;
end process;
process (clock_c) begin
  if rising_edge(clock_c) then
    if i5 = "1" then
      n6 <= "0";
    elsif i4 = "1" then
      n6 <= n5;
    end if;
  end if;
end process;
n7 <= s29_1(10 downto 10) &
  s29_1(9 downto 9) &
  s29_1(8 downto 8) &
  s29_1(7 downto 7) &
  s29_1(6 downto 6) &
  s29_1(5 downto 5) &
  s29_1(4 downto 4) &
  s29_1(3 downto 3) &
  s29_1(2 downto 2) &
  s29_1(1 downto 1);
process (clock_c) begin
  if rising_edge(clock_c) then
    if i5 = "1" then
      n8 <= "0000000000";
    elsif i4 = "1" then
      n8 <= n7;
    end if;
  end if;
end process;
process (clock_c) begin
  if rising_edge(clock_c) then
    if i5 = "1" then
      n9 <= "0000000000";
    elsif i4 = "1" then
      n9 <= n8;
    end if;
  end if;
end process;
process (clock_c) begin
  if rising_edge(clock_c) then
    if i5 = "1" then
      n10 <= "0000000000";
    elsif i4 = "1" then
      n10 <= n9;
    end if;
  end if;
end process;
process (clock_c) begin
  if rising_edge(clock_c) then
    if i5 = "1" then
      n11 <= "0000000000";
    elsif i4 = "1" then
      n11 <= n10;
    end if;
  end if;
end process;
n12 <= s29_1(0 downto 0);
process (clock_c) begin
  if rising_edge(clock_c) then
    if i5 = "1" then
      n13 <= "0";
    elsif i4 = "1" then
      n13 <= n12;
    end if;
  end if;
end process;
process (clock_c) begin
  if rising_edge(clock_c) then
    if i5 = "1" then
      n14 <= "0";
    elsif i4 = "1" then
      n14 <= n13;
    end if;
  end if;
end process;
process (clock_c) begin
  if rising_edge(clock_c) then
    if i5 = "1" then
      n15 <= "0";
    elsif i4 = "1" then
      n15 <= n14;
    end if;
  end if;
end process;
process (clock_c) begin
  if rising_edge(clock_c) then
    if i5 = "1" then
      n16 <= "0";
    elsif i4 = "1" then
      n16 <= n15;
    end if;
  end if;
end process;
n17 <= not n16;
n18 <= s28_2 & s28_1;
n19 <= s28_3(71 downto 71) &
  s28_3(70 downto 70) &
  s28_3(69 downto 69) &
  s28_3(68 downto 68) &
  s28_3(67 downto 67) &
  s28_3(66 downto 66) &
  s28_3(65 downto 65) &
  s28_3(64 downto 64) &
  s28_3(63 downto 63) &
  s28_3(62 downto 62) &
  s28_3(61 downto 61) &
  s28_3(60 downto 60) &
  s28_3(59 downto 59) &
  s28_3(58 downto 58) &
  s28_3(57 downto 57) &
  s28_3(56 downto 56) &
  s28_3(55 downto 55) &
  s28_3(54 downto 54) &
  s28_3(53 downto 53) &
  s28_3(52 downto 52) &
  s28_3(51 downto 51) &
  s28_3(50 downto 50) &
  s28_3(49 downto 49) &
  s28_3(48 downto 48) &
  s28_3(47 downto 47) &
  s28_3(46 downto 46) &
  s28_3(45 downto 45) &
  s28_3(44 downto 44) &
  s28_3(43 downto 43) &
  s28_3(42 downto 42) &
  s28_3(41 downto 41) &
  s28_3(40 downto 40) &
  s28_3(39 downto 39) &
  s28_3(38 downto 38) &
  s28_3(37 downto 37) &
  s28_3(36 downto 36);
n20 <= s28_3(35 downto 35) &
  s28_3(34 downto 34) &
  s28_3(33 downto 33) &
  s28_3(32 downto 32) &
  s28_3(31 downto 31) &
  s28_3(30 downto 30) &
  s28_3(29 downto 29) &
  s28_3(28 downto 28) &
  s28_3(27 downto 27) &
  s28_3(26 downto 26) &
  s28_3(25 downto 25) &
  s28_3(24 downto 24) &
  s28_3(23 downto 23) &
  s28_3(22 downto 22) &
  s28_3(21 downto 21) &
  s28_3(20 downto 20) &
  s28_3(19 downto 19) &
  s28_3(18 downto 18) &
  s28_3(17 downto 17) &
  s28_3(16 downto 16) &
  s28_3(15 downto 15) &
  s28_3(14 downto 14) &
  s28_3(13 downto 13) &
  s28_3(12 downto 12) &
  s28_3(11 downto 11) &
  s28_3(10 downto 10) &
  s28_3(9 downto 9) &
  s28_3(8 downto 8) &
  s28_3(7 downto 7) &
  s28_3(6 downto 6) &
  s28_3(5 downto 5) &
  s28_3(4 downto 4) &
  s28_3(3 downto 3) &
  s28_3(2 downto 2) &
  s28_3(1 downto 1) &
  s28_3(0 downto 0);
n21 <= s27_1(71 downto 71) &
  s27_1(70 downto 70) &
  s27_1(69 downto 69) &
  s27_1(68 downto 68) &
  s27_1(67 downto 67) &
  s27_1(66 downto 66) &
  s27_1(65 downto 65) &
  s27_1(64 downto 64) &
  s27_1(63 downto 63) &
  s27_1(62 downto 62) &
  s27_1(61 downto 61) &
  s27_1(60 downto 60) &
  s27_1(59 downto 59) &
  s27_1(58 downto 58) &
  s27_1(57 downto 57) &
  s27_1(56 downto 56) &
  s27_1(55 downto 55) &
  s27_1(54 downto 54) &
  s27_1(53 downto 53) &
  s27_1(52 downto 52) &
  s27_1(51 downto 51) &
  s27_1(50 downto 50) &
  s27_1(49 downto 49) &
  s27_1(48 downto 48) &
  s27_1(47 downto 47) &
  s27_1(46 downto 46) &
  s27_1(45 downto 45) &
  s27_1(44 downto 44) &
  s27_1(43 downto 43) &
  s27_1(42 downto 42) &
  s27_1(41 downto 41) &
  s27_1(40 downto 40) &
  s27_1(39 downto 39) &
  s27_1(38 downto 38) &
  s27_1(37 downto 37) &
  s27_1(36 downto 36);
n22 <= s27_1(35 downto 35) &
  s27_1(34 downto 34) &
  s27_1(33 downto 33) &
  s27_1(32 downto 32) &
  s27_1(31 downto 31) &
  s27_1(30 downto 30) &
  s27_1(29 downto 29) &
  s27_1(28 downto 28) &
  s27_1(27 downto 27) &
  s27_1(26 downto 26) &
  s27_1(25 downto 25) &
  s27_1(24 downto 24) &
  s27_1(23 downto 23) &
  s27_1(22 downto 22) &
  s27_1(21 downto 21) &
  s27_1(20 downto 20) &
  s27_1(19 downto 19) &
  s27_1(18 downto 18) &
  s27_1(17 downto 17) &
  s27_1(16 downto 16) &
  s27_1(15 downto 15) &
  s27_1(14 downto 14) &
  s27_1(13 downto 13) &
  s27_1(12 downto 12) &
  s27_1(11 downto 11) &
  s27_1(10 downto 10) &
  s27_1(9 downto 9) &
  s27_1(8 downto 8) &
  s27_1(7 downto 7) &
  s27_1(6 downto 6) &
  s27_1(5 downto 5) &
  s27_1(4 downto 4) &
  s27_1(3 downto 3) &
  s27_1(2 downto 2) &
  s27_1(1 downto 1) &
  s27_1(0 downto 0);
n23 <= n20 when s26_1 = "1" else n19;
n24 <= n22 when s26_1 = "1" else n21;
s25 : cf_fft_4096_18_43 port map (clock_c, i2, i3, n1, i4, i5, s25_1, s25_2);
s26 : cf_fft_4096_18_37 port map (clock_c, n18, i4, i5, s26_1);
s27 : cf_fft_4096_18_33 port map (clock_c, n2, n6, n11, n16, i4, i5, s27_1);
s28 : cf_fft_4096_18_32 port map (clock_c, n2, n6, n11, n17, i4, i5, s28_1, s28_2, s28_3);
s29 : cf_fft_4096_18_28 port map (clock_c, i1, i4, i5, s29_1, s29_2);
o3 <= n24;
o2 <= n23;
o1 <= s28_1;
end architecture rtl;

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
entity cf_fft_4096_18_26 is
port (
clock_c : in std_logic;
i1 : in  unsigned(35 downto 0);
i2 : in  unsigned(35 downto 0);
i3 : in  unsigned(10 downto 0);
i4 : in  unsigned(0 downto 0);
i5 : in  unsigned(0 downto 0);
o1 : out unsigned(35 downto 0);
o2 : out unsigned(35 downto 0));
end entity cf_fft_4096_18_26;
architecture rtl of cf_fft_4096_18_26 is
signal n1 : unsigned(35 downto 0) := "000000000000000000000000000000000000";
signal n2 : unsigned(17 downto 0);
signal n3 : unsigned(17 downto 0);
signal n4 : unsigned(35 downto 0) := "000000000000000000000000000000000000";
signal n5 : unsigned(17 downto 0);
signal n6 : unsigned(17 downto 0);
signal n7 : unsigned(17 downto 0) := "000000000000000000";
signal n8 : unsigned(17 downto 0) := "000000000000000000";
signal n9 : unsigned(17 downto 0) := "000000000000000000";
signal n10 : unsigned(17 downto 0) := "000000000000000000";
signal n11 : unsigned(35 downto 0) := "000000000000000000000000000000000000";
signal n12 : unsigned(17 downto 0);
signal n13 : unsigned(17 downto 0);
signal n14 : unsigned(35 downto 0);
signal n15 : unsigned(17 downto 0);
signal n16 : unsigned(17 downto 0) := "000000000000000000";
signal n17 : unsigned(35 downto 0);
signal n18 : unsigned(17 downto 0);
signal n19 : unsigned(17 downto 0) := "000000000000000000";
signal n20 : unsigned(17 downto 0);
signal n21 : unsigned(17 downto 0) := "000000000000000000";
signal n22 : unsigned(35 downto 0);
signal n23 : unsigned(17 downto 0);
signal n24 : unsigned(17 downto 0) := "000000000000000000";
signal n25 : unsigned(35 downto 0);
signal n26 : unsigned(17 downto 0);
signal n27 : unsigned(17 downto 0) := "000000000000000000";
signal n28 : unsigned(17 downto 0);
signal n29 : unsigned(17 downto 0) := "000000000000000000";
signal n30 : unsigned(17 downto 0);
signal n31 : unsigned(17 downto 0);
signal n32 : unsigned(35 downto 0);
signal n33 : unsigned(35 downto 0) := "000000000000000000000000000000000000";
signal n34 : unsigned(17 downto 0);
signal n35 : unsigned(17 downto 0);
signal n36 : unsigned(35 downto 0);
signal n37 : unsigned(35 downto 0) := "000000000000000000000000000000000000";
begin
process (clock_c) begin
  if rising_edge(clock_c) then
    if i5 = "1" then
      n1 <= "000000000000000000000000000000000000";
    elsif i4 = "1" then
      n1 <= i1;
    end if;
  end if;
end process;
n2 <= n1(35 downto 35) &
  n1(34 downto 34) &
  n1(33 downto 33) &
  n1(32 downto 32) &
  n1(31 downto 31) &
  n1(30 downto 30) &
  n1(29 downto 29) &
  n1(28 downto 28) &
  n1(27 downto 27) &
  n1(26 downto 26) &
  n1(25 downto 25) &
  n1(24 downto 24) &
  n1(23 downto 23) &
  n1(22 downto 22) &
  n1(21 downto 21) &
  n1(20 downto 20) &
  n1(19 downto 19) &
  n1(18 downto 18);
n3 <= n1(17 downto 17) &
  n1(16 downto 16) &
  n1(15 downto 15) &
  n1(14 downto 14) &
  n1(13 downto 13) &
  n1(12 downto 12) &
  n1(11 downto 11) &
  n1(10 downto 10) &
  n1(9 downto 9) &
  n1(8 downto 8) &
  n1(7 downto 7) &
  n1(6 downto 6) &
  n1(5 downto 5) &
  n1(4 downto 4) &
  n1(3 downto 3) &
  n1(2 downto 2) &
  n1(1 downto 1) &
  n1(0 downto 0);
process (clock_c) begin
  if rising_edge(clock_c) then
    if i5 = "1" then
      n4 <= "000000000000000000000000000000000000";
    elsif i4 = "1" then
      n4 <= i2;
    end if;
  end if;
end process;
n5 <= n4(35 downto 35) &
  n4(34 downto 34) &
  n4(33 downto 33) &
  n4(32 downto 32) &
  n4(31 downto 31) &
  n4(30 downto 30) &
  n4(29 downto 29) &
  n4(28 downto 28) &
  n4(27 downto 27) &
  n4(26 downto 26) &
  n4(25 downto 25) &
  n4(24 downto 24) &
  n4(23 downto 23) &
  n4(22 downto 22) &
  n4(21 downto 21) &
  n4(20 downto 20) &
  n4(19 downto 19) &
  n4(18 downto 18);
n6 <= n4(17 downto 17) &
  n4(16 downto 16) &
  n4(15 downto 15) &
  n4(14 downto 14) &
  n4(13 downto 13) &
  n4(12 downto 12) &
  n4(11 downto 11) &
  n4(10 downto 10) &
  n4(9 downto 9) &
  n4(8 downto 8) &
  n4(7 downto 7) &
  n4(6 downto 6) &
  n4(5 downto 5) &
  n4(4 downto 4) &
  n4(3 downto 3) &
  n4(2 downto 2) &
  n4(1 downto 1) &
  n4(0 downto 0);
process (clock_c) begin
  if rising_edge(clock_c) then
    if i5 = "1" then
      n7 <= "000000000000000000";
    elsif i4 = "1" then
      n7 <= n2;
    end if;
  end if;
end process;
process (clock_c) begin
  if rising_edge(clock_c) then
    if i5 = "1" then
      n8 <= "000000000000000000";
    elsif i4 = "1" then
      n8 <= n7;
    end if;
  end if;
end process;
process (clock_c) begin
  if rising_edge(clock_c) then
    if i5 = "1" then
      n9 <= "000000000000000000";
    elsif i4 = "1" then
      n9 <= n3;
    end if;
  end if;
end process;
process (clock_c) begin
  if rising_edge(clock_c) then
    if i5 = "1" then
      n10 <= "000000000000000000";
    elsif i4 = "1" then
      n10 <= n9;
    end if;
  end if;
end process;
process (clock_c) begin
  if rising_edge(clock_c) then 
    if i4 = "1" then
      case i3 is
        when "00000000000" => n11 <= "011111111111111111000000000000000000";
        when "00000000001" => n11 <= "011111111111111111111111111100110110";
        when "00000000010" => n11 <= "011111111111111111111111111001101101";
        when "00000000011" => n11 <= "011111111111111110111111110110100100";
        when "00000000100" => n11 <= "011111111111111101111111110011011011";
        when "00000000101" => n11 <= "011111111111111100111111110000010010";
        when "00000000110" => n11 <= "011111111111111010111111101101001001";
        when "00000000111" => n11 <= "011111111111111000111111101010000000";
        when "00000001000" => n11 <= "011111111111110110111111100110110111";
        when "00000001001" => n11 <= "011111111111110011111111100011101110";
        when "00000001010" => n11 <= "011111111111110000111111100000100101";
        when "00000001011" => n11 <= "011111111111101101111111011101011100";
        when "00000001100" => n11 <= "011111111111101001111111011010010011";
        when "00000001101" => n11 <= "011111111111100101111111010111001010";
        when "00000001110" => n11 <= "011111111111100001111111010100000001";
        when "00000001111" => n11 <= "011111111111011101111111010000111000";
        when "00000010000" => n11 <= "011111111111011000111111001101101111";
        when "00000010001" => n11 <= "011111111111010011111111001010100110";
        when "00000010010" => n11 <= "011111111111001110111111000111011101";
        when "00000010011" => n11 <= "011111111111001000111111000100010100";
        when "00000010100" => n11 <= "011111111111000010111111000001001011";
        when "00000010101" => n11 <= "011111111110111011111110111110000010";
        when "00000010110" => n11 <= "011111111110110101111110111010111001";
        when "00000010111" => n11 <= "011111111110101110111110110111110000";
        when "00000011000" => n11 <= "011111111110100111111110110100100111";
        when "00000011001" => n11 <= "011111111110011111111110110001011110";
        when "00000011010" => n11 <= "011111111110010111111110101110010101";
        when "00000011011" => n11 <= "011111111110001111111110101011001100";
        when "00000011100" => n11 <= "011111111110000111111110101000000011";
        when "00000011101" => n11 <= "011111111101111110111110100100111011";
        when "00000011110" => n11 <= "011111111101110101111110100001110010";
        when "00000011111" => n11 <= "011111111101101011111110011110101001";
        when "00000100000" => n11 <= "011111111101100010111110011011100000";
        when "00000100001" => n11 <= "011111111101011000111110011000010111";
        when "00000100010" => n11 <= "011111111101001101111110010101001110";
        when "00000100011" => n11 <= "011111111101000011111110010010000110";
        when "00000100100" => n11 <= "011111111100111000111110001110111101";
        when "00000100101" => n11 <= "011111111100101100111110001011110100";
        when "00000100110" => n11 <= "011111111100100001111110001000101011";
        when "00000100111" => n11 <= "011111111100010101111110000101100011";
        when "00000101000" => n11 <= "011111111100001001111110000010011010";
        when "00000101001" => n11 <= "011111111011111100111101111111010001";
        when "00000101010" => n11 <= "011111111011110000111101111100001001";
        when "00000101011" => n11 <= "011111111011100010111101111001000000";
        when "00000101100" => n11 <= "011111111011010101111101110101110111";
        when "00000101101" => n11 <= "011111111011000111111101110010101111";
        when "00000101110" => n11 <= "011111111010111001111101101111100110";
        when "00000101111" => n11 <= "011111111010101011111101101100011110";
        when "00000110000" => n11 <= "011111111010011100111101101001010101";
        when "00000110001" => n11 <= "011111111010001101111101100110001101";
        when "00000110010" => n11 <= "011111111001111110111101100011000100";
        when "00000110011" => n11 <= "011111111001101111111101011111111100";
        when "00000110100" => n11 <= "011111111001011111111101011100110011";
        when "00000110101" => n11 <= "011111111001001111111101011001101011";
        when "00000110110" => n11 <= "011111111000111110111101010110100011";
        when "00000110111" => n11 <= "011111111000101101111101010011011010";
        when "00000111000" => n11 <= "011111111000011100111101010000010010";
        when "00000111001" => n11 <= "011111111000001011111101001101001010";
        when "00000111010" => n11 <= "011111110111111001111101001010000001";
        when "00000111011" => n11 <= "011111110111100111111101000110111001";
        when "00000111100" => n11 <= "011111110111010101111101000011110001";
        when "00000111101" => n11 <= "011111110111000010111101000000101001";
        when "00000111110" => n11 <= "011111110110101111111100111101100000";
        when "00000111111" => n11 <= "011111110110011100111100111010011000";
        when "00001000000" => n11 <= "011111110110001000111100110111010000";
        when "00001000001" => n11 <= "011111110101110100111100110100001000";
        when "00001000010" => n11 <= "011111110101100000111100110001000000";
        when "00001000011" => n11 <= "011111110101001100111100101101111000";
        when "00001000100" => n11 <= "011111110100110111111100101010110000";
        when "00001000101" => n11 <= "011111110100100010111100100111101000";
        when "00001000110" => n11 <= "011111110100001101111100100100100000";
        when "00001000111" => n11 <= "011111110011110111111100100001011000";
        when "00001001000" => n11 <= "011111110011100001111100011110010000";
        when "00001001001" => n11 <= "011111110011001011111100011011001001";
        when "00001001010" => n11 <= "011111110010110100111100011000000001";
        when "00001001011" => n11 <= "011111110010011101111100010100111001";
        when "00001001100" => n11 <= "011111110010000110111100010001110001";
        when "00001001101" => n11 <= "011111110001101110111100001110101010";
        when "00001001110" => n11 <= "011111110001010110111100001011100010";
        when "00001001111" => n11 <= "011111110000111110111100001000011010";
        when "00001010000" => n11 <= "011111110000100110111100000101010011";
        when "00001010001" => n11 <= "011111110000001101111100000010001011";
        when "00001010010" => n11 <= "011111101111110100111011111111000100";
        when "00001010011" => n11 <= "011111101111011011111011111011111100";
        when "00001010100" => n11 <= "011111101111000001111011111000110101";
        when "00001010101" => n11 <= "011111101110100111111011110101101110";
        when "00001010110" => n11 <= "011111101110001101111011110010100110";
        when "00001010111" => n11 <= "011111101101110010111011101111011111";
        when "00001011000" => n11 <= "011111101101010111111011101100011000";
        when "00001011001" => n11 <= "011111101100111100111011101001010001";
        when "00001011010" => n11 <= "011111101100100000111011100110001001";
        when "00001011011" => n11 <= "011111101100000101111011100011000010";
        when "00001011100" => n11 <= "011111101011101000111011011111111011";
        when "00001011101" => n11 <= "011111101011001100111011011100110100";
        when "00001011110" => n11 <= "011111101010101111111011011001101101";
        when "00001011111" => n11 <= "011111101010010010111011010110100110";
        when "00001100000" => n11 <= "011111101001110101111011010011011111";
        when "00001100001" => n11 <= "011111101001010111111011010000011000";
        when "00001100010" => n11 <= "011111101000111001111011001101010010";
        when "00001100011" => n11 <= "011111101000011011111011001010001011";
        when "00001100100" => n11 <= "011111100111111100111011000111000100";
        when "00001100101" => n11 <= "011111100111011110111011000011111101";
        when "00001100110" => n11 <= "011111100110111110111011000000110111";
        when "00001100111" => n11 <= "011111100110011111111010111101110000";
        when "00001101000" => n11 <= "011111100101111111111010111010101010";
        when "00001101001" => n11 <= "011111100101011111111010110111100011";
        when "00001101010" => n11 <= "011111100100111111111010110100011101";
        when "00001101011" => n11 <= "011111100100011110111010110001010110";
        when "00001101100" => n11 <= "011111100011111101111010101110010000";
        when "00001101101" => n11 <= "011111100011011100111010101011001010";
        when "00001101110" => n11 <= "011111100010111010111010101000000011";
        when "00001101111" => n11 <= "011111100010011000111010100100111101";
        when "00001110000" => n11 <= "011111100001110110111010100001110111";
        when "00001110001" => n11 <= "011111100001010011111010011110110001";
        when "00001110010" => n11 <= "011111100000110000111010011011101011";
        when "00001110011" => n11 <= "011111100000001101111010011000100101";
        when "00001110100" => n11 <= "011111011111101010111010010101011111";
        when "00001110101" => n11 <= "011111011111000110111010010010011001";
        when "00001110110" => n11 <= "011111011110100010111010001111010100";
        when "00001110111" => n11 <= "011111011101111110111010001100001110";
        when "00001111000" => n11 <= "011111011101011001111010001001001000";
        when "00001111001" => n11 <= "011111011100110100111010000110000010";
        when "00001111010" => n11 <= "011111011100001111111010000010111101";
        when "00001111011" => n11 <= "011111011011101001111001111111110111";
        when "00001111100" => n11 <= "011111011011000011111001111100110010";
        when "00001111101" => n11 <= "011111011010011101111001111001101100";
        when "00001111110" => n11 <= "011111011001110111111001110110100111";
        when "00001111111" => n11 <= "011111011001010000111001110011100010";
        when "00010000000" => n11 <= "011111011000101001111001110000011101";
        when "00010000001" => n11 <= "011111011000000010111001101101010111";
        when "00010000010" => n11 <= "011111010111011010111001101010010010";
        when "00010000011" => n11 <= "011111010110110010111001100111001101";
        when "00010000100" => n11 <= "011111010110001010111001100100001000";
        when "00010000101" => n11 <= "011111010101100001111001100001000011";
        when "00010000110" => n11 <= "011111010100111000111001011101111111";
        when "00010000111" => n11 <= "011111010100001111111001011010111010";
        when "00010001000" => n11 <= "011111010011100110111001010111110101";
        when "00010001001" => n11 <= "011111010010111100111001010100110000";
        when "00010001010" => n11 <= "011111010010010010111001010001101100";
        when "00010001011" => n11 <= "011111010001100111111001001110100111";
        when "00010001100" => n11 <= "011111010000111101111001001011100011";
        when "00010001101" => n11 <= "011111010000010010111001001000011110";
        when "00010001110" => n11 <= "011111001111100110111001000101011010";
        when "00010001111" => n11 <= "011111001110111011111001000010010110";
        when "00010010000" => n11 <= "011111001110001111111000111111010001";
        when "00010010001" => n11 <= "011111001101100011111000111100001101";
        when "00010010010" => n11 <= "011111001100110110111000111001001001";
        when "00010010011" => n11 <= "011111001100001001111000110110000101";
        when "00010010100" => n11 <= "011111001011011100111000110011000001";
        when "00010010101" => n11 <= "011111001010101111111000101111111101";
        when "00010010110" => n11 <= "011111001010000001111000101100111010";
        when "00010010111" => n11 <= "011111001001010011111000101001110110";
        when "00010011000" => n11 <= "011111001000100101111000100110110010";
        when "00010011001" => n11 <= "011111000111110110111000100011101111";
        when "00010011010" => n11 <= "011111000111000111111000100000101011";
        when "00010011011" => n11 <= "011111000110011000111000011101101000";
        when "00010011100" => n11 <= "011111000101101000111000011010100100";
        when "00010011101" => n11 <= "011111000100111001111000010111100001";
        when "00010011110" => n11 <= "011111000100001001111000010100011110";
        when "00010011111" => n11 <= "011111000011011000111000010001011011";
        when "00010100000" => n11 <= "011111000010100111111000001110011000";
        when "00010100001" => n11 <= "011111000001110110111000001011010101";
        when "00010100010" => n11 <= "011111000001000101111000001000010010";
        when "00010100011" => n11 <= "011111000000010100111000000101001111";
        when "00010100100" => n11 <= "011110111111100010111000000010001100";
        when "00010100101" => n11 <= "011110111110101111110111111111001001";
        when "00010100110" => n11 <= "011110111101111101110111111100000111";
        when "00010100111" => n11 <= "011110111101001010110111111001000100";
        when "00010101000" => n11 <= "011110111100010111110111110110000010";
        when "00010101001" => n11 <= "011110111011100100110111110010111111";
        when "00010101010" => n11 <= "011110111010110000110111101111111101";
        when "00010101011" => n11 <= "011110111001111100110111101100111011";
        when "00010101100" => n11 <= "011110111001001000110111101001111001";
        when "00010101101" => n11 <= "011110111000010011110111100110110111";
        when "00010101110" => n11 <= "011110110111011110110111100011110101";
        when "00010101111" => n11 <= "011110110110101001110111100000110011";
        when "00010110000" => n11 <= "011110110101110100110111011101110001";
        when "00010110001" => n11 <= "011110110100111110110111011010101111";
        when "00010110010" => n11 <= "011110110100001000110111010111101110";
        when "00010110011" => n11 <= "011110110011010001110111010100101100";
        when "00010110100" => n11 <= "011110110010011011110111010001101010";
        when "00010110101" => n11 <= "011110110001100100110111001110101001";
        when "00010110110" => n11 <= "011110110000101100110111001011101000";
        when "00010110111" => n11 <= "011110101111110101110111001000100111";
        when "00010111000" => n11 <= "011110101110111101110111000101100101";
        when "00010111001" => n11 <= "011110101110000101110111000010100100";
        when "00010111010" => n11 <= "011110101101001100110110111111100011";
        when "00010111011" => n11 <= "011110101100010100110110111100100010";
        when "00010111100" => n11 <= "011110101011011011110110111001100010";
        when "00010111101" => n11 <= "011110101010100001110110110110100001";
        when "00010111110" => n11 <= "011110101001101000110110110011100000";
        when "00010111111" => n11 <= "011110101000101110110110110000100000";
        when "00011000000" => n11 <= "011110100111110100110110101101011111";
        when "00011000001" => n11 <= "011110100110111001110110101010011111";
        when "00011000010" => n11 <= "011110100101111110110110100111011111";
        when "00011000011" => n11 <= "011110100101000011110110100100011110";
        when "00011000100" => n11 <= "011110100100001000110110100001011110";
        when "00011000101" => n11 <= "011110100011001100110110011110011110";
        when "00011000110" => n11 <= "011110100010010000110110011011011111";
        when "00011000111" => n11 <= "011110100001010100110110011000011111";
        when "00011001000" => n11 <= "011110100000010111110110010101011111";
        when "00011001001" => n11 <= "011110011111011010110110010010011111";
        when "00011001010" => n11 <= "011110011110011101110110001111100000";
        when "00011001011" => n11 <= "011110011101100000110110001100100000";
        when "00011001100" => n11 <= "011110011100100010110110001001100001";
        when "00011001101" => n11 <= "011110011011100100110110000110100010";
        when "00011001110" => n11 <= "011110011010100110110110000011100011";
        when "00011001111" => n11 <= "011110011001100111110110000000100100";
        when "00011010000" => n11 <= "011110011000101000110101111101100101";
        when "00011010001" => n11 <= "011110010111101001110101111010100110";
        when "00011010010" => n11 <= "011110010110101001110101110111100111";
        when "00011010011" => n11 <= "011110010101101010110101110100101000";
        when "00011010100" => n11 <= "011110010100101001110101110001101010";
        when "00011010101" => n11 <= "011110010011101001110101101110101011";
        when "00011010110" => n11 <= "011110010010101000110101101011101101";
        when "00011010111" => n11 <= "011110010001100111110101101000101111";
        when "00011011000" => n11 <= "011110010000100110110101100101110000";
        when "00011011001" => n11 <= "011110001111100101110101100010110010";
        when "00011011010" => n11 <= "011110001110100011110101011111110100";
        when "00011011011" => n11 <= "011110001101100001110101011100110111";
        when "00011011100" => n11 <= "011110001100011110110101011001111001";
        when "00011011101" => n11 <= "011110001011011011110101010110111011";
        when "00011011110" => n11 <= "011110001010011000110101010011111101";
        when "00011011111" => n11 <= "011110001001010101110101010001000000";
        when "00011100000" => n11 <= "011110001000010010110101001110000011";
        when "00011100001" => n11 <= "011110000111001110110101001011000101";
        when "00011100010" => n11 <= "011110000110001010110101001000001000";
        when "00011100011" => n11 <= "011110000101000101110101000101001011";
        when "00011100100" => n11 <= "011110000100000000110101000010001110";
        when "00011100101" => n11 <= "011110000010111011110100111111010001";
        when "00011100110" => n11 <= "011110000001110110110100111100010101";
        when "00011100111" => n11 <= "011110000000110000110100111001011000";
        when "00011101000" => n11 <= "011101111111101010110100110110011100";
        when "00011101001" => n11 <= "011101111110100100110100110011011111";
        when "00011101010" => n11 <= "011101111101011110110100110000100011";
        when "00011101011" => n11 <= "011101111100010111110100101101100111";
        when "00011101100" => n11 <= "011101111011010000110100101010101011";
        when "00011101101" => n11 <= "011101111010001001110100100111101111";
        when "00011101110" => n11 <= "011101111001000001110100100100110011";
        when "00011101111" => n11 <= "011101110111111001110100100001110111";
        when "00011110000" => n11 <= "011101110110110001110100011110111011";
        when "00011110001" => n11 <= "011101110101101000110100011100000000";
        when "00011110010" => n11 <= "011101110100011111110100011001000100";
        when "00011110011" => n11 <= "011101110011010110110100010110001001";
        when "00011110100" => n11 <= "011101110010001101110100010011001110";
        when "00011110101" => n11 <= "011101110001000011110100010000010011";
        when "00011110110" => n11 <= "011101101111111001110100001101011000";
        when "00011110111" => n11 <= "011101101110101111110100001010011101";
        when "00011111000" => n11 <= "011101101101100101110100000111100010";
        when "00011111001" => n11 <= "011101101100011010110100000100101000";
        when "00011111010" => n11 <= "011101101011001111110100000001101101";
        when "00011111011" => n11 <= "011101101010000011110011111110110011";
        when "00011111100" => n11 <= "011101101000111000110011111011111000";
        when "00011111101" => n11 <= "011101100111101100110011111000111110";
        when "00011111110" => n11 <= "011101100110100000110011110110000100";
        when "00011111111" => n11 <= "011101100101010011110011110011001010";
        when "00100000000" => n11 <= "011101100100000110110011110000010000";
        when "00100000001" => n11 <= "011101100010111001110011101101010111";
        when "00100000010" => n11 <= "011101100001101100110011101010011101";
        when "00100000011" => n11 <= "011101100000011110110011100111100100";
        when "00100000100" => n11 <= "011101011111010000110011100100101010";
        when "00100000101" => n11 <= "011101011110000010110011100001110001";
        when "00100000110" => n11 <= "011101011100110011110011011110111000";
        when "00100000111" => n11 <= "011101011011100101110011011011111111";
        when "00100001000" => n11 <= "011101011010010110110011011001000110";
        when "00100001001" => n11 <= "011101011001000110110011010110001101";
        when "00100001010" => n11 <= "011101010111110111110011010011010101";
        when "00100001011" => n11 <= "011101010110100111110011010000011100";
        when "00100001100" => n11 <= "011101010101010110110011001101100100";
        when "00100001101" => n11 <= "011101010100000110110011001010101100";
        when "00100001110" => n11 <= "011101010010110101110011000111110100";
        when "00100001111" => n11 <= "011101010001100100110011000100111100";
        when "00100010000" => n11 <= "011101010000010011110011000010000100";
        when "00100010001" => n11 <= "011101001111000001110010111111001100";
        when "00100010010" => n11 <= "011101001101101111110010111100010100";
        when "00100010011" => n11 <= "011101001100011101110010111001011101";
        when "00100010100" => n11 <= "011101001011001011110010110110100101";
        when "00100010101" => n11 <= "011101001001111000110010110011101110";
        when "00100010110" => n11 <= "011101001000100101110010110000110111";
        when "00100010111" => n11 <= "011101000111010010110010101110000000";
        when "00100011000" => n11 <= "011101000101111110110010101011001001";
        when "00100011001" => n11 <= "011101000100101010110010101000010011";
        when "00100011010" => n11 <= "011101000011010110110010100101011100";
        when "00100011011" => n11 <= "011101000010000010110010100010100101";
        when "00100011100" => n11 <= "011101000000101101110010011111101111";
        when "00100011101" => n11 <= "011100111111011000110010011100111001";
        when "00100011110" => n11 <= "011100111110000011110010011010000011";
        when "00100011111" => n11 <= "011100111100101101110010010111001101";
        when "00100100000" => n11 <= "011100111011010111110010010100010111";
        when "00100100001" => n11 <= "011100111010000001110010010001100001";
        when "00100100010" => n11 <= "011100111000101011110010001110101100";
        when "00100100011" => n11 <= "011100110111010100110010001011110110";
        when "00100100100" => n11 <= "011100110101111101110010001001000001";
        when "00100100101" => n11 <= "011100110100100110110010000110001100";
        when "00100100110" => n11 <= "011100110011001110110010000011010111";
        when "00100100111" => n11 <= "011100110001110111110010000000100010";
        when "00100101000" => n11 <= "011100110000011111110001111101101101";
        when "00100101001" => n11 <= "011100101111000110110001111010111001";
        when "00100101010" => n11 <= "011100101101101110110001111000000100";
        when "00100101011" => n11 <= "011100101100010101110001110101010000";
        when "00100101100" => n11 <= "011100101010111100110001110010011100";
        when "00100101101" => n11 <= "011100101001100010110001101111100111";
        when "00100101110" => n11 <= "011100101000001000110001101100110100";
        when "00100101111" => n11 <= "011100100110101110110001101010000000";
        when "00100110000" => n11 <= "011100100101010100110001100111001100";
        when "00100110001" => n11 <= "011100100011111010110001100100011001";
        when "00100110010" => n11 <= "011100100010011111110001100001100101";
        when "00100110011" => n11 <= "011100100001000100110001011110110010";
        when "00100110100" => n11 <= "011100011111101000110001011011111111";
        when "00100110101" => n11 <= "011100011110001101110001011001001100";
        when "00100110110" => n11 <= "011100011100110001110001010110011001";
        when "00100110111" => n11 <= "011100011011010101110001010011100110";
        when "00100111000" => n11 <= "011100011001111000110001010000110100";
        when "00100111001" => n11 <= "011100011000011011110001001110000001";
        when "00100111010" => n11 <= "011100010110111110110001001011001111";
        when "00100111011" => n11 <= "011100010101100001110001001000011101";
        when "00100111100" => n11 <= "011100010100000100110001000101101011";
        when "00100111101" => n11 <= "011100010010100110110001000010111001";
        when "00100111110" => n11 <= "011100010001001000110001000000001000";
        when "00100111111" => n11 <= "011100001111101001110000111101010110";
        when "00101000000" => n11 <= "011100001110001011110000111010100101";
        when "00101000001" => n11 <= "011100001100101100110000110111110011";
        when "00101000010" => n11 <= "011100001011001101110000110101000010";
        when "00101000011" => n11 <= "011100001001101101110000110010010001";
        when "00101000100" => n11 <= "011100001000001101110000101111100000";
        when "00101000101" => n11 <= "011100000110101101110000101100110000";
        when "00101000110" => n11 <= "011100000101001101110000101001111111";
        when "00101000111" => n11 <= "011100000011101101110000100111001111";
        when "00101001000" => n11 <= "011100000010001100110000100100011111";
        when "00101001001" => n11 <= "011100000000101011110000100001101111";
        when "00101001010" => n11 <= "011011111111001001110000011110111111";
        when "00101001011" => n11 <= "011011111101101000110000011100001111";
        when "00101001100" => n11 <= "011011111100000110110000011001011111";
        when "00101001101" => n11 <= "011011111010100100110000010110110000";
        when "00101001110" => n11 <= "011011111001000001110000010100000001";
        when "00101001111" => n11 <= "011011110111011111110000010001010001";
        when "00101010000" => n11 <= "011011110101111100110000001110100010";
        when "00101010001" => n11 <= "011011110100011000110000001011110011";
        when "00101010010" => n11 <= "011011110010110101110000001001000101";
        when "00101010011" => n11 <= "011011110001010001110000000110010110";
        when "00101010100" => n11 <= "011011101111101101110000000011101000";
        when "00101010101" => n11 <= "011011101110001001110000000000111010";
        when "00101010110" => n11 <= "011011101100100100101111111110001011";
        when "00101010111" => n11 <= "011011101010111111101111111011011110";
        when "00101011000" => n11 <= "011011101001011010101111111000110000";
        when "00101011001" => n11 <= "011011100111110101101111110110000010";
        when "00101011010" => n11 <= "011011100110001111101111110011010101";
        when "00101011011" => n11 <= "011011100100101001101111110000100111";
        when "00101011100" => n11 <= "011011100011000011101111101101111010";
        when "00101011101" => n11 <= "011011100001011101101111101011001101";
        when "00101011110" => n11 <= "011011011111110110101111101000100000";
        when "00101011111" => n11 <= "011011011110001111101111100101110100";
        when "00101100000" => n11 <= "011011011100101000101111100011000111";
        when "00101100001" => n11 <= "011011011011000000101111100000011011";
        when "00101100010" => n11 <= "011011011001011000101111011101101110";
        when "00101100011" => n11 <= "011011010111110000101111011011000010";
        when "00101100100" => n11 <= "011011010110001000101111011000010110";
        when "00101100101" => n11 <= "011011010100100000101111010101101011";
        when "00101100110" => n11 <= "011011010010110111101111010010111111";
        when "00101100111" => n11 <= "011011010001001110101111010000010100";
        when "00101101000" => n11 <= "011011001111100100101111001101101000";
        when "00101101001" => n11 <= "011011001101111011101111001010111101";
        when "00101101010" => n11 <= "011011001100010001101111001000010010";
        when "00101101011" => n11 <= "011011001010100111101111000101101000";
        when "00101101100" => n11 <= "011011001000111100101111000010111101";
        when "00101101101" => n11 <= "011011000111010010101111000000010011";
        when "00101101110" => n11 <= "011011000101100111101110111101101000";
        when "00101101111" => n11 <= "011011000011111100101110111010111110";
        when "00101110000" => n11 <= "011011000010010000101110111000010100";
        when "00101110001" => n11 <= "011011000000100100101110110101101011";
        when "00101110010" => n11 <= "011010111110111000101110110011000001";
        when "00101110011" => n11 <= "011010111101001100101110110000010111";
        when "00101110100" => n11 <= "011010111011100000101110101101101110";
        when "00101110101" => n11 <= "011010111001110011101110101011000101";
        when "00101110110" => n11 <= "011010111000000110101110101000011100";
        when "00101110111" => n11 <= "011010110110011001101110100101110011";
        when "00101111000" => n11 <= "011010110100101011101110100011001011";
        when "00101111001" => n11 <= "011010110010111110101110100000100010";
        when "00101111010" => n11 <= "011010110001001111101110011101111010";
        when "00101111011" => n11 <= "011010101111100001101110011011010010";
        when "00101111100" => n11 <= "011010101101110011101110011000101010";
        when "00101111101" => n11 <= "011010101100000100101110010110000010";
        when "00101111110" => n11 <= "011010101010010101101110010011011010";
        when "00101111111" => n11 <= "011010101000100101101110010000110011";
        when "00110000000" => n11 <= "011010100110110110101110001110001100";
        when "00110000001" => n11 <= "011010100101000110101110001011100101";
        when "00110000010" => n11 <= "011010100011010110101110001000111110";
        when "00110000011" => n11 <= "011010100001100110101110000110010111";
        when "00110000100" => n11 <= "011010011111110101101110000011110000";
        when "00110000101" => n11 <= "011010011110000100101110000001001010";
        when "00110000110" => n11 <= "011010011100010011101101111110100100";
        when "00110000111" => n11 <= "011010011010100010101101111011111110";
        when "00110001000" => n11 <= "011010011000110000101101111001011000";
        when "00110001001" => n11 <= "011010010110111110101101110110110010";
        when "00110001010" => n11 <= "011010010101001100101101110100001101";
        when "00110001011" => n11 <= "011010010011011010101101110001100111";
        when "00110001100" => n11 <= "011010010001100111101101101111000010";
        when "00110001101" => n11 <= "011010001111110100101101101100011101";
        when "00110001110" => n11 <= "011010001110000001101101101001111000";
        when "00110001111" => n11 <= "011010001100001110101101100111010100";
        when "00110010000" => n11 <= "011010001010011010101101100100101111";
        when "00110010001" => n11 <= "011010001000100110101101100010001011";
        when "00110010010" => n11 <= "011010000110110010101101011111100111";
        when "00110010011" => n11 <= "011010000100111110101101011101000011";
        when "00110010100" => n11 <= "011010000011001001101101011010011111";
        when "00110010101" => n11 <= "011010000001010100101101010111111011";
        when "00110010110" => n11 <= "011001111111011111101101010101011000";
        when "00110010111" => n11 <= "011001111101101001101101010010110101";
        when "00110011000" => n11 <= "011001111011110100101101010000010010";
        when "00110011001" => n11 <= "011001111001111110101101001101101111";
        when "00110011010" => n11 <= "011001111000001000101101001011001100";
        when "00110011011" => n11 <= "011001110110010001101101001000101010";
        when "00110011100" => n11 <= "011001110100011011101101000110000111";
        when "00110011101" => n11 <= "011001110010100100101101000011100101";
        when "00110011110" => n11 <= "011001110000101101101101000001000011";
        when "00110011111" => n11 <= "011001101110110101101100111110100010";
        when "00110100000" => n11 <= "011001101100111110101100111100000000";
        when "00110100001" => n11 <= "011001101011000110101100111001011111";
        when "00110100010" => n11 <= "011001101001001101101100110110111101";
        when "00110100011" => n11 <= "011001100111010101101100110100011100";
        when "00110100100" => n11 <= "011001100101011100101100110001111011";
        when "00110100101" => n11 <= "011001100011100100101100101111011011";
        when "00110100110" => n11 <= "011001100001101010101100101100111010";
        when "00110100111" => n11 <= "011001011111110001101100101010011010";
        when "00110101000" => n11 <= "011001011101110111101100100111111010";
        when "00110101001" => n11 <= "011001011011111110101100100101011010";
        when "00110101010" => n11 <= "011001011010000011101100100010111010";
        when "00110101011" => n11 <= "011001011000001001101100100000011011";
        when "00110101100" => n11 <= "011001010110001110101100011101111011";
        when "00110101101" => n11 <= "011001010100010100101100011011011100";
        when "00110101110" => n11 <= "011001010010011001101100011000111101";
        when "00110101111" => n11 <= "011001010000011101101100010110011110";
        when "00110110000" => n11 <= "011001001110100010101100010100000000";
        when "00110110001" => n11 <= "011001001100100110101100010001100001";
        when "00110110010" => n11 <= "011001001010101010101100001111000011";
        when "00110110011" => n11 <= "011001001000101101101100001100100101";
        when "00110110100" => n11 <= "011001000110110001101100001010000111";
        when "00110110101" => n11 <= "011001000100110100101100000111101010";
        when "00110110110" => n11 <= "011001000010110111101100000101001100";
        when "00110110111" => n11 <= "011001000000111010101100000010101111";
        when "00110111000" => n11 <= "011000111110111100101100000000010010";
        when "00110111001" => n11 <= "011000111100111111101011111101110101";
        when "00110111010" => n11 <= "011000111011000001101011111011011000";
        when "00110111011" => n11 <= "011000111001000010101011111000111100";
        when "00110111100" => n11 <= "011000110111000100101011110110100000";
        when "00110111101" => n11 <= "011000110101000101101011110100000011";
        when "00110111110" => n11 <= "011000110011000110101011110001101000";
        when "00110111111" => n11 <= "011000110001000111101011101111001100";
        when "00111000000" => n11 <= "011000101111001000101011101100110000";
        when "00111000001" => n11 <= "011000101101001000101011101010010101";
        when "00111000010" => n11 <= "011000101011001000101011100111111010";
        when "00111000011" => n11 <= "011000101001001000101011100101011111";
        when "00111000100" => n11 <= "011000100111000111101011100011000100";
        when "00111000101" => n11 <= "011000100101000111101011100000101010";
        when "00111000110" => n11 <= "011000100011000110101011011110001111";
        when "00111000111" => n11 <= "011000100001000101101011011011110101";
        when "00111001000" => n11 <= "011000011111000100101011011001011011";
        when "00111001001" => n11 <= "011000011101000010101011010111000001";
        when "00111001010" => n11 <= "011000011011000000101011010100101000";
        when "00111001011" => n11 <= "011000011000111110101011010010001111";
        when "00111001100" => n11 <= "011000010110111100101011001111110101";
        when "00111001101" => n11 <= "011000010100111001101011001101011100";
        when "00111001110" => n11 <= "011000010010110111101011001011000100";
        when "00111001111" => n11 <= "011000010000110100101011001000101011";
        when "00111010000" => n11 <= "011000001110110000101011000110010011";
        when "00111010001" => n11 <= "011000001100101101101011000011111011";
        when "00111010010" => n11 <= "011000001010101001101011000001100011";
        when "00111010011" => n11 <= "011000001000100101101010111111001011";
        when "00111010100" => n11 <= "011000000110100001101010111100110011";
        when "00111010101" => n11 <= "011000000100011101101010111010011100";
        when "00111010110" => n11 <= "011000000010011000101010111000000101";
        when "00111010111" => n11 <= "011000000000010011101010110101101110";
        when "00111011000" => n11 <= "010111111110001110101010110011010111";
        when "00111011001" => n11 <= "010111111100001001101010110001000001";
        when "00111011010" => n11 <= "010111111010000011101010101110101011";
        when "00111011011" => n11 <= "010111110111111110101010101100010100";
        when "00111011100" => n11 <= "010111110101111000101010101001111110";
        when "00111011101" => n11 <= "010111110011110001101010100111101001";
        when "00111011110" => n11 <= "010111110001101011101010100101010011";
        when "00111011111" => n11 <= "010111101111100100101010100010111110";
        when "00111100000" => n11 <= "010111101101011101101010100000101001";
        when "00111100001" => n11 <= "010111101011010110101010011110010100";
        when "00111100010" => n11 <= "010111101001001111101010011011111111";
        when "00111100011" => n11 <= "010111100111000111101010011001101011";
        when "00111100100" => n11 <= "010111100101000000101010010111010111";
        when "00111100101" => n11 <= "010111100010110111101010010101000011";
        when "00111100110" => n11 <= "010111100000101111101010010010101111";
        when "00111100111" => n11 <= "010111011110100111101010010000011011";
        when "00111101000" => n11 <= "010111011100011110101010001110001000";
        when "00111101001" => n11 <= "010111011010010101101010001011110101";
        when "00111101010" => n11 <= "010111011000001100101010001001100010";
        when "00111101011" => n11 <= "010111010110000010101010000111001111";
        when "00111101100" => n11 <= "010111010011111001101010000100111100";
        when "00111101101" => n11 <= "010111010001101111101010000010101010";
        when "00111101110" => n11 <= "010111001111100101101010000000011000";
        when "00111101111" => n11 <= "010111001101011011101001111110000110";
        when "00111110000" => n11 <= "010111001011010000101001111011110100";
        when "00111110001" => n11 <= "010111001001000101101001111001100011";
        when "00111110010" => n11 <= "010111000110111010101001110111010001";
        when "00111110011" => n11 <= "010111000100101111101001110101000000";
        when "00111110100" => n11 <= "010111000010100100101001110010101111";
        when "00111110101" => n11 <= "010111000000011000101001110000011111";
        when "00111110110" => n11 <= "010110111110001100101001101110001110";
        when "00111110111" => n11 <= "010110111100000000101001101011111110";
        when "00111111000" => n11 <= "010110111001110100101001101001101110";
        when "00111111001" => n11 <= "010110110111100111101001100111011110";
        when "00111111010" => n11 <= "010110110101011010101001100101001111";
        when "00111111011" => n11 <= "010110110011001110101001100010111111";
        when "00111111100" => n11 <= "010110110001000000101001100000110000";
        when "00111111101" => n11 <= "010110101110110011101001011110100001";
        when "00111111110" => n11 <= "010110101100100101101001011100010010";
        when "00111111111" => n11 <= "010110101010010111101001011010000100";
        when "01000000000" => n11 <= "010110101000001001101001010111110110";
        when "01000000001" => n11 <= "010110100101111011101001010101101000";
        when "01000000010" => n11 <= "010110100011101101101001010011011010";
        when "01000000011" => n11 <= "010110100001011110101001010001001100";
        when "01000000100" => n11 <= "010110011111001111101001001110111111";
        when "01000000101" => n11 <= "010110011101000000101001001100110001";
        when "01000000110" => n11 <= "010110011010110000101001001010100101";
        when "01000000111" => n11 <= "010110011000100001101001001000011000";
        when "01000001000" => n11 <= "010110010110010001101001000110001011";
        when "01000001001" => n11 <= "010110010100000001101001000011111111";
        when "01000001010" => n11 <= "010110010001110001101001000001110011";
        when "01000001011" => n11 <= "010110001111100000101000111111100111";
        when "01000001100" => n11 <= "010110001101010000101000111101011011";
        when "01000001101" => n11 <= "010110001010111111101000111011010000";
        when "01000001110" => n11 <= "010110001000101110101000111001000101";
        when "01000001111" => n11 <= "010110000110011100101000110110111010";
        when "01000010000" => n11 <= "010110000100001011101000110100101111";
        when "01000010001" => n11 <= "010110000001111001101000110010100100";
        when "01000010010" => n11 <= "010101111111100111101000110000011010";
        when "01000010011" => n11 <= "010101111101010101101000101110010000";
        when "01000010100" => n11 <= "010101111011000011101000101100000110";
        when "01000010101" => n11 <= "010101111000110000101000101001111101";
        when "01000010110" => n11 <= "010101110110011101101000100111110011";
        when "01000010111" => n11 <= "010101110100001010101000100101101010";
        when "01000011000" => n11 <= "010101110001110111101000100011100001";
        when "01000011001" => n11 <= "010101101111100100101000100001011000";
        when "01000011010" => n11 <= "010101101101010000101000011111010000";
        when "01000011011" => n11 <= "010101101010111100101000011101001000";
        when "01000011100" => n11 <= "010101101000101000101000011010111111";
        when "01000011101" => n11 <= "010101100110010100101000011000111000";
        when "01000011110" => n11 <= "010101100100000000101000010110110000";
        when "01000011111" => n11 <= "010101100001101011101000010100101001";
        when "01000100000" => n11 <= "010101011111010110101000010010100010";
        when "01000100001" => n11 <= "010101011101000001101000010000011011";
        when "01000100010" => n11 <= "010101011010101100101000001110010100";
        when "01000100011" => n11 <= "010101011000010110101000001100001110";
        when "01000100100" => n11 <= "010101010110000001101000001010000111";
        when "01000100101" => n11 <= "010101010011101011101000001000000001";
        when "01000100110" => n11 <= "010101010001010100101000000101111100";
        when "01000100111" => n11 <= "010101001110111110101000000011110110";
        when "01000101000" => n11 <= "010101001100101000101000000001110001";
        when "01000101001" => n11 <= "010101001010010001100111111111101100";
        when "01000101010" => n11 <= "010101000111111010100111111101100111";
        when "01000101011" => n11 <= "010101000101100011100111111011100010";
        when "01000101100" => n11 <= "010101000011001100100111111001011110";
        when "01000101101" => n11 <= "010101000000110100100111110111011010";
        when "01000101110" => n11 <= "010100111110011100100111110101010110";
        when "01000101111" => n11 <= "010100111100000100100111110011010010";
        when "01000110000" => n11 <= "010100111001101100100111110001001111";
        when "01000110001" => n11 <= "010100110111010100100111101111001011";
        when "01000110010" => n11 <= "010100110100111011100111101101001000";
        when "01000110011" => n11 <= "010100110010100011100111101011000110";
        when "01000110100" => n11 <= "010100110000001010100111101001000011";
        when "01000110101" => n11 <= "010100101101110000100111100111000001";
        when "01000110110" => n11 <= "010100101011010111100111100100111111";
        when "01000110111" => n11 <= "010100101000111110100111100010111101";
        when "01000111000" => n11 <= "010100100110100100100111100000111011";
        when "01000111001" => n11 <= "010100100100001010100111011110111010";
        when "01000111010" => n11 <= "010100100001110000100111011100111001";
        when "01000111011" => n11 <= "010100011111010101100111011010111000";
        when "01000111100" => n11 <= "010100011100111011100111011000111000";
        when "01000111101" => n11 <= "010100011010100000100111010110110111";
        when "01000111110" => n11 <= "010100011000000101100111010100110111";
        when "01000111111" => n11 <= "010100010101101010100111010010110111";
        when "01001000000" => n11 <= "010100010011001111100111010000110111";
        when "01001000001" => n11 <= "010100010000110011100111001110111000";
        when "01001000010" => n11 <= "010100001110010111100111001100111001";
        when "01001000011" => n11 <= "010100001011111100100111001010111010";
        when "01001000100" => n11 <= "010100001001011111100111001000111011";
        when "01001000101" => n11 <= "010100000111000011100111000110111101";
        when "01001000110" => n11 <= "010100000100100111100111000100111110";
        when "01001000111" => n11 <= "010100000010001010100111000011000000";
        when "01001001000" => n11 <= "010011111111101101100111000001000011";
        when "01001001001" => n11 <= "010011111101010000100110111111000101";
        when "01001001010" => n11 <= "010011111010110011100110111101001000";
        when "01001001011" => n11 <= "010011111000010101100110111011001011";
        when "01001001100" => n11 <= "010011110101111000100110111001001110";
        when "01001001101" => n11 <= "010011110011011010100110110111010010";
        when "01001001110" => n11 <= "010011110000111100100110110101010101";
        when "01001001111" => n11 <= "010011101110011110100110110011011001";
        when "01001010000" => n11 <= "010011101011111111100110110001011101";
        when "01001010001" => n11 <= "010011101001100001100110101111100010";
        when "01001010010" => n11 <= "010011100111000010100110101101100110";
        when "01001010011" => n11 <= "010011100100100011100110101011101011";
        when "01001010100" => n11 <= "010011100010000100100110101001110001";
        when "01001010101" => n11 <= "010011011111100100100110100111110110";
        when "01001010110" => n11 <= "010011011101000101100110100101111100";
        when "01001010111" => n11 <= "010011011010100101100110100100000001";
        when "01001011000" => n11 <= "010011011000000101100110100010001000";
        when "01001011001" => n11 <= "010011010101100101100110100000001110";
        when "01001011010" => n11 <= "010011010011000101100110011110010101";
        when "01001011011" => n11 <= "010011010000100100100110011100011011";
        when "01001011100" => n11 <= "010011001110000100100110011010100011";
        when "01001011101" => n11 <= "010011001011100011100110011000101010";
        when "01001011110" => n11 <= "010011001001000010100110010110110010";
        when "01001011111" => n11 <= "010011000110100000100110010100111001";
        when "01001100000" => n11 <= "010011000011111111100110010011000001";
        when "01001100001" => n11 <= "010011000001011101100110010001001010";
        when "01001100010" => n11 <= "010010111110111100100110001111010010";
        when "01001100011" => n11 <= "010010111100011010100110001101011011";
        when "01001100100" => n11 <= "010010111001111000100110001011100100";
        when "01001100101" => n11 <= "010010110111010101100110001001101110";
        when "01001100110" => n11 <= "010010110100110011100110000111110111";
        when "01001100111" => n11 <= "010010110010010000100110000110000001";
        when "01001101000" => n11 <= "010010101111101101100110000100001011";
        when "01001101001" => n11 <= "010010101101001010100110000010010110";
        when "01001101010" => n11 <= "010010101010100111100110000000100000";
        when "01001101011" => n11 <= "010010101000000100100101111110101011";
        when "01001101100" => n11 <= "010010100101100000100101111100110110";
        when "01001101101" => n11 <= "010010100010111100100101111011000001";
        when "01001101110" => n11 <= "010010100000011000100101111001001101";
        when "01001101111" => n11 <= "010010011101110100100101110111011001";
        when "01001110000" => n11 <= "010010011011010000100101110101100101";
        when "01001110001" => n11 <= "010010011000101011100101110011110001";
        when "01001110010" => n11 <= "010010010110000111100101110001111110";
        when "01001110011" => n11 <= "010010010011100010100101110000001011";
        when "01001110100" => n11 <= "010010010000111101100101101110011000";
        when "01001110101" => n11 <= "010010001110011000100101101100100101";
        when "01001110110" => n11 <= "010010001011110010100101101010110011";
        when "01001110111" => n11 <= "010010001001001101100101101001000001";
        when "01001111000" => n11 <= "010010000110100111100101100111001111";
        when "01001111001" => n11 <= "010010000100000001100101100101011101";
        when "01001111010" => n11 <= "010010000001011011100101100011101100";
        when "01001111011" => n11 <= "010001111110110101100101100001111011";
        when "01001111100" => n11 <= "010001111100001111100101100000001010";
        when "01001111101" => n11 <= "010001111001101000100101011110011001";
        when "01001111110" => n11 <= "010001110111000001100101011100101001";
        when "01001111111" => n11 <= "010001110100011010100101011010111001";
        when "01010000000" => n11 <= "010001110001110011100101011001001001";
        when "01010000001" => n11 <= "010001101111001100100101010111011010";
        when "01010000010" => n11 <= "010001101100100101100101010101101010";
        when "01010000011" => n11 <= "010001101001111101100101010011111011";
        when "01010000100" => n11 <= "010001100111010101100101010010001100";
        when "01010000101" => n11 <= "010001100100101101100101010000011110";
        when "01010000110" => n11 <= "010001100010000101100101001110110000";
        when "01010000111" => n11 <= "010001011111011101100101001101000001";
        when "01010001000" => n11 <= "010001011100110100100101001011010100";
        when "01010001001" => n11 <= "010001011010001100100101001001100110";
        when "01010001010" => n11 <= "010001010111100011100101000111111001";
        when "01010001011" => n11 <= "010001010100111010100101000110001100";
        when "01010001100" => n11 <= "010001010010010001100101000100011111";
        when "01010001101" => n11 <= "010001001111101000100101000010110011";
        when "01010001110" => n11 <= "010001001100111110100101000001000111";
        when "01010001111" => n11 <= "010001001010010100100100111111011011";
        when "01010010000" => n11 <= "010001000111101011100100111101101111";
        when "01010010001" => n11 <= "010001000101000001100100111100000011";
        when "01010010010" => n11 <= "010001000010010111100100111010011000";
        when "01010010011" => n11 <= "010000111111101100100100111000101101";
        when "01010010100" => n11 <= "010000111101000010100100110111000011";
        when "01010010101" => n11 <= "010000111010010111100100110101011000";
        when "01010010110" => n11 <= "010000110111101101100100110011101110";
        when "01010010111" => n11 <= "010000110101000010100100110010000100";
        when "01010011000" => n11 <= "010000110010010111100100110000011011";
        when "01010011001" => n11 <= "010000101111101011100100101110110001";
        when "01010011010" => n11 <= "010000101101000000100100101101001000";
        when "01010011011" => n11 <= "010000101010010100100100101011011111";
        when "01010011100" => n11 <= "010000100111101001100100101001110111";
        when "01010011101" => n11 <= "010000100100111101100100101000001111";
        when "01010011110" => n11 <= "010000100010010001100100100110100111";
        when "01010011111" => n11 <= "010000011111100100100100100100111111";
        when "01010100000" => n11 <= "010000011100111000100100100011010111";
        when "01010100001" => n11 <= "010000011010001011100100100001110000";
        when "01010100010" => n11 <= "010000010111011111100100100000001001";
        when "01010100011" => n11 <= "010000010100110010100100011110100010";
        when "01010100100" => n11 <= "010000010010000101100100011100111100";
        when "01010100101" => n11 <= "010000001111011000100100011011010110";
        when "01010100110" => n11 <= "010000001100101010100100011001110000";
        when "01010100111" => n11 <= "010000001001111101100100011000001010";
        when "01010101000" => n11 <= "010000000111001111100100010110100101";
        when "01010101001" => n11 <= "010000000100100001100100010101000000";
        when "01010101010" => n11 <= "010000000001110100100100010011011011";
        when "01010101011" => n11 <= "001111111111000101100100010001110110";
        when "01010101100" => n11 <= "001111111100010111100100010000010010";
        when "01010101101" => n11 <= "001111111001101001100100001110101110";
        when "01010101110" => n11 <= "001111110110111010100100001101001010";
        when "01010101111" => n11 <= "001111110100001100100100001011100111";
        when "01010110000" => n11 <= "001111110001011101100100001010000011";
        when "01010110001" => n11 <= "001111101110101110100100001000100000";
        when "01010110010" => n11 <= "001111101011111110100100000110111110";
        when "01010110011" => n11 <= "001111101001001111100100000101011011";
        when "01010110100" => n11 <= "001111100110100000100100000011111001";
        when "01010110101" => n11 <= "001111100011110000100100000010010111";
        when "01010110110" => n11 <= "001111100001000000100100000000110110";
        when "01010110111" => n11 <= "001111011110010000100011111111010100";
        when "01010111000" => n11 <= "001111011011100000100011111101110011";
        when "01010111001" => n11 <= "001111011000110000100011111100010010";
        when "01010111010" => n11 <= "001111010110000000100011111010110010";
        when "01010111011" => n11 <= "001111010011001111100011111001010010";
        when "01010111100" => n11 <= "001111010000011111100011110111110010";
        when "01010111101" => n11 <= "001111001101101110100011110110010010";
        when "01010111110" => n11 <= "001111001010111101100011110100110010";
        when "01010111111" => n11 <= "001111001000001100100011110011010011";
        when "01011000000" => n11 <= "001111000101011010100011110001110100";
        when "01011000001" => n11 <= "001111000010101001100011110000010110";
        when "01011000010" => n11 <= "001110111111110111100011101110110111";
        when "01011000011" => n11 <= "001110111101000110100011101101011001";
        when "01011000100" => n11 <= "001110111010010100100011101011111011";
        when "01011000101" => n11 <= "001110110111100010100011101010011110";
        when "01011000110" => n11 <= "001110110100110000100011101001000001";
        when "01011000111" => n11 <= "001110110001111110100011100111100100";
        when "01011001000" => n11 <= "001110101111001011100011100110000111";
        when "01011001001" => n11 <= "001110101100011001100011100100101010";
        when "01011001010" => n11 <= "001110101001100110100011100011001110";
        when "01011001011" => n11 <= "001110100110110011100011100001110010";
        when "01011001100" => n11 <= "001110100100000000100011100000010111";
        when "01011001101" => n11 <= "001110100001001101100011011110111011";
        when "01011001110" => n11 <= "001110011110011010100011011101100000";
        when "01011001111" => n11 <= "001110011011100110100011011100000101";
        when "01011010000" => n11 <= "001110011000110011100011011010101011";
        when "01011010001" => n11 <= "001110010101111111100011011001010001";
        when "01011010010" => n11 <= "001110010011001011100011010111110111";
        when "01011010011" => n11 <= "001110010000011000100011010110011101";
        when "01011010100" => n11 <= "001110001101100011100011010101000011";
        when "01011010101" => n11 <= "001110001010101111100011010011101010";
        when "01011010110" => n11 <= "001110000111111011100011010010010001";
        when "01011010111" => n11 <= "001110000101000110100011010000111001";
        when "01011011000" => n11 <= "001110000010010010100011001111100000";
        when "01011011001" => n11 <= "001101111111011101100011001110001000";
        when "01011011010" => n11 <= "001101111100101000100011001100110001";
        when "01011011011" => n11 <= "001101111001110011100011001011011001";
        when "01011011100" => n11 <= "001101110110111110100011001010000010";
        when "01011011101" => n11 <= "001101110100001001100011001000101011";
        when "01011011110" => n11 <= "001101110001010011100011000111010100";
        when "01011011111" => n11 <= "001101101110011110100011000101111110";
        when "01011100000" => n11 <= "001101101011101000100011000100101000";
        when "01011100001" => n11 <= "001101101000110010100011000011010010";
        when "01011100010" => n11 <= "001101100101111100100011000001111100";
        when "01011100011" => n11 <= "001101100011000110100011000000100111";
        when "01011100100" => n11 <= "001101100000010000100010111111010010";
        when "01011100101" => n11 <= "001101011101011010100010111101111101";
        when "01011100110" => n11 <= "001101011010100011100010111100101001";
        when "01011100111" => n11 <= "001101010111101100100010111011010101";
        when "01011101000" => n11 <= "001101010100110110100010111010000001";
        when "01011101001" => n11 <= "001101010001111111100010111000101101";
        when "01011101010" => n11 <= "001101001111001000100010110111011010";
        when "01011101011" => n11 <= "001101001100010001100010110110000111";
        when "01011101100" => n11 <= "001101001001011010100010110100110100";
        when "01011101101" => n11 <= "001101000110100010100010110011100010";
        when "01011101110" => n11 <= "001101000011101011100010110010010000";
        when "01011101111" => n11 <= "001101000000110011100010110000111110";
        when "01011110000" => n11 <= "001100111101111011100010101111101100";
        when "01011110001" => n11 <= "001100111011000011100010101110011011";
        when "01011110010" => n11 <= "001100111000001011100010101101001010";
        when "01011110011" => n11 <= "001100110101010011100010101011111001";
        when "01011110100" => n11 <= "001100110010011011100010101010101001";
        when "01011110101" => n11 <= "001100101111100011100010101001011000";
        when "01011110110" => n11 <= "001100101100101010100010101000001000";
        when "01011110111" => n11 <= "001100101001110010100010100110111001";
        when "01011111000" => n11 <= "001100100110111001100010100101101001";
        when "01011111001" => n11 <= "001100100100000000100010100100011010";
        when "01011111010" => n11 <= "001100100001000111100010100011001100";
        when "01011111011" => n11 <= "001100011110001110100010100001111101";
        when "01011111100" => n11 <= "001100011011010101100010100000101111";
        when "01011111101" => n11 <= "001100011000011011100010011111100001";
        when "01011111110" => n11 <= "001100010101100010100010011110010011";
        when "01011111111" => n11 <= "001100010010101000100010011101000110";
        when "01100000000" => n11 <= "001100001111101111100010011011111001";
        when "01100000001" => n11 <= "001100001100110101100010011010101100";
        when "01100000010" => n11 <= "001100001001111011100010011001011111";
        when "01100000011" => n11 <= "001100000111000001100010011000010011";
        when "01100000100" => n11 <= "001100000100000111100010010111000111";
        when "01100000101" => n11 <= "001100000001001100100010010101111100";
        when "01100000110" => n11 <= "001011111110010010100010010100110000";
        when "01100000111" => n11 <= "001011111011010111100010010011100101";
        when "01100001000" => n11 <= "001011111000011101100010010010011010";
        when "01100001001" => n11 <= "001011110101100010100010010001010000";
        when "01100001010" => n11 <= "001011110010100111100010010000000110";
        when "01100001011" => n11 <= "001011101111101100100010001110111100";
        when "01100001100" => n11 <= "001011101100110001100010001101110010";
        when "01100001101" => n11 <= "001011101001110110100010001100101001";
        when "01100001110" => n11 <= "001011100110111011100010001011100000";
        when "01100001111" => n11 <= "001011100011111111100010001010010111";
        when "01100010000" => n11 <= "001011100001000100100010001001001110";
        when "01100010001" => n11 <= "001011011110001000100010001000000110";
        when "01100010010" => n11 <= "001011011011001100100010000110111110";
        when "01100010011" => n11 <= "001011011000010000100010000101110110";
        when "01100010100" => n11 <= "001011010101010100100010000100101111";
        when "01100010101" => n11 <= "001011010010011000100010000011101000";
        when "01100010110" => n11 <= "001011001111011100100010000010100001";
        when "01100010111" => n11 <= "001011001100100000100010000001011011";
        when "01100011000" => n11 <= "001011001001100011100010000000010101";
        when "01100011001" => n11 <= "001011000110100111100001111111001111";
        when "01100011010" => n11 <= "001011000011101010100001111110001001";
        when "01100011011" => n11 <= "001011000000101110100001111101000100";
        when "01100011100" => n11 <= "001010111101110001100001111011111111";
        when "01100011101" => n11 <= "001010111010110100100001111010111010";
        when "01100011110" => n11 <= "001010110111110111100001111001110101";
        when "01100011111" => n11 <= "001010110100111010100001111000110001";
        when "01100100000" => n11 <= "001010110001111100100001110111101101";
        when "01100100001" => n11 <= "001010101110111111100001110110101010";
        when "01100100010" => n11 <= "001010101100000010100001110101100111";
        when "01100100011" => n11 <= "001010101001000100100001110100100100";
        when "01100100100" => n11 <= "001010100110000110100001110011100001";
        when "01100100101" => n11 <= "001010100011001000100001110010011110";
        when "01100100110" => n11 <= "001010100000001011100001110001011100";
        when "01100100111" => n11 <= "001010011101001101100001110000011010";
        when "01100101000" => n11 <= "001010011010001111100001101111011001";
        when "01100101001" => n11 <= "001010010111010000100001101110011000";
        when "01100101010" => n11 <= "001010010100010010100001101101010111";
        when "01100101011" => n11 <= "001010010001010100100001101100010110";
        when "01100101100" => n11 <= "001010001110010101100001101011010110";
        when "01100101101" => n11 <= "001010001011010111100001101010010101";
        when "01100101110" => n11 <= "001010001000011000100001101001010110";
        when "01100101111" => n11 <= "001010000101011001100001101000010110";
        when "01100110000" => n11 <= "001010000010011010100001100111010111";
        when "01100110001" => n11 <= "001001111111011011100001100110011000";
        when "01100110010" => n11 <= "001001111100011100100001100101011001";
        when "01100110011" => n11 <= "001001111001011101100001100100011011";
        when "01100110100" => n11 <= "001001110110011110100001100011011101";
        when "01100110101" => n11 <= "001001110011011111100001100010011111";
        when "01100110110" => n11 <= "001001110000011111100001100001100010";
        when "01100110111" => n11 <= "001001101101100000100001100000100101";
        when "01100111000" => n11 <= "001001101010100000100001011111101000";
        when "01100111001" => n11 <= "001001100111100000100001011110101011";
        when "01100111010" => n11 <= "001001100100100000100001011101101111";
        when "01100111011" => n11 <= "001001100001100001100001011100110011";
        when "01100111100" => n11 <= "001001011110100001100001011011110111";
        when "01100111101" => n11 <= "001001011011100001100001011010111100";
        when "01100111110" => n11 <= "001001011000100000100001011010000001";
        when "01100111111" => n11 <= "001001010101100000100001011001000110";
        when "01101000000" => n11 <= "001001010010100000100001011000001011";
        when "01101000001" => n11 <= "001001001111011111100001010111010001";
        when "01101000010" => n11 <= "001001001100011111100001010110010111";
        when "01101000011" => n11 <= "001001001001011110100001010101011110";
        when "01101000100" => n11 <= "001001000110011101100001010100100100";
        when "01101000101" => n11 <= "001001000011011101100001010011101011";
        when "01101000110" => n11 <= "001001000000011100100001010010110011";
        when "01101000111" => n11 <= "001000111101011011100001010001111010";
        when "01101001000" => n11 <= "001000111010011010100001010001000010";
        when "01101001001" => n11 <= "001000110111011000100001010000001010";
        when "01101001010" => n11 <= "001000110100010111100001001111010011";
        when "01101001011" => n11 <= "001000110001010110100001001110011011";
        when "01101001100" => n11 <= "001000101110010101100001001101100100";
        when "01101001101" => n11 <= "001000101011010011100001001100101110";
        when "01101001110" => n11 <= "001000101000010001100001001011110111";
        when "01101001111" => n11 <= "001000100101010000100001001011000001";
        when "01101010000" => n11 <= "001000100010001110100001001010001011";
        when "01101010001" => n11 <= "001000011111001100100001001001010110";
        when "01101010010" => n11 <= "001000011100001010100001001000100001";
        when "01101010011" => n11 <= "001000011001001000100001000111101100";
        when "01101010100" => n11 <= "001000010110000110100001000110110111";
        when "01101010101" => n11 <= "001000010011000100100001000110000011";
        when "01101010110" => n11 <= "001000010000000010100001000101001111";
        when "01101010111" => n11 <= "001000001101000000100001000100011011";
        when "01101011000" => n11 <= "001000001001111101100001000011101000";
        when "01101011001" => n11 <= "001000000110111011100001000010110101";
        when "01101011010" => n11 <= "001000000011111000100001000010000010";
        when "01101011011" => n11 <= "001000000000110110100001000001010000";
        when "01101011100" => n11 <= "000111111101110011100001000000011101";
        when "01101011101" => n11 <= "000111111010110000100000111111101011";
        when "01101011110" => n11 <= "000111110111101101100000111110111010";
        when "01101011111" => n11 <= "000111110100101010100000111110001001";
        when "01101100000" => n11 <= "000111110001100111100000111101011000";
        when "01101100001" => n11 <= "000111101110100100100000111100100111";
        when "01101100010" => n11 <= "000111101011100001100000111011110110";
        when "01101100011" => n11 <= "000111101000011110100000111011000110";
        when "01101100100" => n11 <= "000111100101011011100000111010010111";
        when "01101100101" => n11 <= "000111100010010111100000111001100111";
        when "01101100110" => n11 <= "000111011111010100100000111000111000";
        when "01101100111" => n11 <= "000111011100010000100000111000001001";
        when "01101101000" => n11 <= "000111011001001101100000110111011010";
        when "01101101001" => n11 <= "000111010110001001100000110110101100";
        when "01101101010" => n11 <= "000111010011000101100000110101111110";
        when "01101101011" => n11 <= "000111010000000010100000110101010000";
        when "01101101100" => n11 <= "000111001100111110100000110100100011";
        when "01101101101" => n11 <= "000111001001111010100000110011110110";
        when "01101101110" => n11 <= "000111000110110110100000110011001001";
        when "01101101111" => n11 <= "000111000011110010100000110010011100";
        when "01101110000" => n11 <= "000111000000101110100000110001110000";
        when "01101110001" => n11 <= "000110111101101001100000110001000100";
        when "01101110010" => n11 <= "000110111010100101100000110000011001";
        when "01101110011" => n11 <= "000110110111100001100000101111101101";
        when "01101110100" => n11 <= "000110110100011100100000101111000010";
        when "01101110101" => n11 <= "000110110001011000100000101110011000";
        when "01101110110" => n11 <= "000110101110010011100000101101101101";
        when "01101110111" => n11 <= "000110101011001111100000101101000011";
        when "01101111000" => n11 <= "000110101000001010100000101100011001";
        when "01101111001" => n11 <= "000110100101000101100000101011110000";
        when "01101111010" => n11 <= "000110100010000000100000101011000111";
        when "01101111011" => n11 <= "000110011110111100100000101010011110";
        when "01101111100" => n11 <= "000110011011110111100000101001110101";
        when "01101111101" => n11 <= "000110011000110010100000101001001101";
        when "01101111110" => n11 <= "000110010101101101100000101000100101";
        when "01101111111" => n11 <= "000110010010101000100000100111111101";
        when "01110000000" => n11 <= "000110001111100010100000100111010110";
        when "01110000001" => n11 <= "000110001100011101100000100110101111";
        when "01110000010" => n11 <= "000110001001011000100000100110001000";
        when "01110000011" => n11 <= "000110000110010011100000100101100010";
        when "01110000100" => n11 <= "000110000011001101100000100100111100";
        when "01110000101" => n11 <= "000110000000001000100000100100010110";
        when "01110000110" => n11 <= "000101111101000010100000100011110000";
        when "01110000111" => n11 <= "000101111001111101100000100011001011";
        when "01110001000" => n11 <= "000101110110110111100000100010100110";
        when "01110001001" => n11 <= "000101110011110001100000100010000001";
        when "01110001010" => n11 <= "000101110000101011100000100001011101";
        when "01110001011" => n11 <= "000101101101100110100000100000111001";
        when "01110001100" => n11 <= "000101101010100000100000100000010101";
        when "01110001101" => n11 <= "000101100111011010100000011111110010";
        when "01110001110" => n11 <= "000101100100010100100000011111001111";
        when "01110001111" => n11 <= "000101100001001110100000011110101100";
        when "01110010000" => n11 <= "000101011110001000100000011110001001";
        when "01110010001" => n11 <= "000101011011000010100000011101100111";
        when "01110010010" => n11 <= "000101010111111100100000011101000101";
        when "01110010011" => n11 <= "000101010100110101100000011100100011";
        when "01110010100" => n11 <= "000101010001101111100000011100000010";
        when "01110010101" => n11 <= "000101001110101001100000011011100001";
        when "01110010110" => n11 <= "000101001011100010100000011011000000";
        when "01110010111" => n11 <= "000101001000011100100000011010100000";
        when "01110011000" => n11 <= "000101000101010101100000011010000000";
        when "01110011001" => n11 <= "000101000010001111100000011001100000";
        when "01110011010" => n11 <= "000100111111001000100000011001000001";
        when "01110011011" => n11 <= "000100111100000010100000011000100001";
        when "01110011100" => n11 <= "000100111000111011100000011000000011";
        when "01110011101" => n11 <= "000100110101110100100000010111100100";
        when "01110011110" => n11 <= "000100110010101101100000010111000110";
        when "01110011111" => n11 <= "000100101111100111100000010110101000";
        when "01110100000" => n11 <= "000100101100100000100000010110001010";
        when "01110100001" => n11 <= "000100101001011001100000010101101101";
        when "01110100010" => n11 <= "000100100110010010100000010101010000";
        when "01110100011" => n11 <= "000100100011001011100000010100110011";
        when "01110100100" => n11 <= "000100100000000100100000010100010111";
        when "01110100101" => n11 <= "000100011100111101100000010011111010";
        when "01110100110" => n11 <= "000100011001110110100000010011011111";
        when "01110100111" => n11 <= "000100010110101110100000010011000011";
        when "01110101000" => n11 <= "000100010011100111100000010010101000";
        when "01110101001" => n11 <= "000100010000100000100000010010001101";
        when "01110101010" => n11 <= "000100001101011001100000010001110010";
        when "01110101011" => n11 <= "000100001010010001100000010001011000";
        when "01110101100" => n11 <= "000100000111001010100000010000111110";
        when "01110101101" => n11 <= "000100000100000011100000010000100100";
        when "01110101110" => n11 <= "000100000000111011100000010000001011";
        when "01110101111" => n11 <= "000011111101110100100000001111110010";
        when "01110110000" => n11 <= "000011111010101100100000001111011001";
        when "01110110001" => n11 <= "000011110111100101100000001111000001";
        when "01110110010" => n11 <= "000011110100011101100000001110101001";
        when "01110110011" => n11 <= "000011110001010101100000001110010001";
        when "01110110100" => n11 <= "000011101110001110100000001101111001";
        when "01110110101" => n11 <= "000011101011000110100000001101100010";
        when "01110110110" => n11 <= "000011100111111110100000001101001011";
        when "01110110111" => n11 <= "000011100100110110100000001100110100";
        when "01110111000" => n11 <= "000011100001101111100000001100011110";
        when "01110111001" => n11 <= "000011011110100111100000001100001000";
        when "01110111010" => n11 <= "000011011011011111100000001011110010";
        when "01110111011" => n11 <= "000011011000010111100000001011011101";
        when "01110111100" => n11 <= "000011010101001111100000001011001000";
        when "01110111101" => n11 <= "000011010010000111100000001010110011";
        when "01110111110" => n11 <= "000011001110111111100000001010011111";
        when "01110111111" => n11 <= "000011001011110111100000001010001011";
        when "01111000000" => n11 <= "000011001000101111100000001001110111";
        when "01111000001" => n11 <= "000011000101100111100000001001100011";
        when "01111000010" => n11 <= "000011000010011111100000001001010000";
        when "01111000011" => n11 <= "000010111111010110100000001000111101";
        when "01111000100" => n11 <= "000010111100001110100000001000101010";
        when "01111000101" => n11 <= "000010111001000110100000001000011000";
        when "01111000110" => n11 <= "000010110101111110100000001000000110";
        when "01111000111" => n11 <= "000010110010110101100000000111110100";
        when "01111001000" => n11 <= "000010101111101101100000000111100011";
        when "01111001001" => n11 <= "000010101100100101100000000111010010";
        when "01111001010" => n11 <= "000010101001011100100000000111000001";
        when "01111001011" => n11 <= "000010100110010100100000000110110000";
        when "01111001100" => n11 <= "000010100011001100100000000110100000";
        when "01111001101" => n11 <= "000010100000000011100000000110010000";
        when "01111001110" => n11 <= "000010011100111011100000000110000001";
        when "01111001111" => n11 <= "000010011001110010100000000101110010";
        when "01111010000" => n11 <= "000010010110101010100000000101100011";
        when "01111010001" => n11 <= "000010010011100001100000000101010100";
        when "01111010010" => n11 <= "000010010000011001100000000101000110";
        when "01111010011" => n11 <= "000010001101010000100000000100111000";
        when "01111010100" => n11 <= "000010001010001000100000000100101010";
        when "01111010101" => n11 <= "000010000110111111100000000100011101";
        when "01111010110" => n11 <= "000010000011110110100000000100001111";
        when "01111010111" => n11 <= "000010000000101110100000000100000011";
        when "01111011000" => n11 <= "000001111101100101100000000011110110";
        when "01111011001" => n11 <= "000001111010011100100000000011101010";
        when "01111011010" => n11 <= "000001110111010100100000000011011110";
        when "01111011011" => n11 <= "000001110100001011100000000011010011";
        when "01111011100" => n11 <= "000001110001000010100000000011000111";
        when "01111011101" => n11 <= "000001101101111001100000000010111100";
        when "01111011110" => n11 <= "000001101010110001100000000010110010";
        when "01111011111" => n11 <= "000001100111101000100000000010100111";
        when "01111100000" => n11 <= "000001100100011111100000000010011101";
        when "01111100001" => n11 <= "000001100001010110100000000010010100";
        when "01111100010" => n11 <= "000001011110001101100000000010001010";
        when "01111100011" => n11 <= "000001011011000100100000000010000001";
        when "01111100100" => n11 <= "000001010111111100100000000001111000";
        when "01111100101" => n11 <= "000001010100110011100000000001110000";
        when "01111100110" => n11 <= "000001010001101010100000000001101000";
        when "01111100111" => n11 <= "000001001110100001100000000001100000";
        when "01111101000" => n11 <= "000001001011011000100000000001011000";
        when "01111101001" => n11 <= "000001001000001111100000000001010001";
        when "01111101010" => n11 <= "000001000101000110100000000001001010";
        when "01111101011" => n11 <= "000001000001111101100000000001000100";
        when "01111101100" => n11 <= "000000111110110100100000000000111101";
        when "01111101101" => n11 <= "000000111011101011100000000000110111";
        when "01111101110" => n11 <= "000000111000100010100000000000110001";
        when "01111101111" => n11 <= "000000110101011001100000000000101100";
        when "01111110000" => n11 <= "000000110010010000100000000000100111";
        when "01111110001" => n11 <= "000000101111000111100000000000100010";
        when "01111110010" => n11 <= "000000101011111110100000000000011110";
        when "01111110011" => n11 <= "000000101000110101100000000000011010";
        when "01111110100" => n11 <= "000000100101101100100000000000010110";
        when "01111110101" => n11 <= "000000100010100011100000000000010010";
        when "01111110110" => n11 <= "000000011111011010100000000000001111";
        when "01111110111" => n11 <= "000000011100010001100000000000001100";
        when "01111111000" => n11 <= "000000011001001000100000000000001001";
        when "01111111001" => n11 <= "000000010101111111100000000000000111";
        when "01111111010" => n11 <= "000000010010110110100000000000000101";
        when "01111111011" => n11 <= "000000001111101101100000000000000011";
        when "01111111100" => n11 <= "000000001100100100100000000000000010";
        when "01111111101" => n11 <= "000000001001011011100000000000000001";
        when "01111111110" => n11 <= "000000000110010010100000000000000000";
        when "01111111111" => n11 <= "000000000011001001100000000000000000";
        when "10000000000" => n11 <= "000000000000000000100000000000000000";
        when "10000000001" => n11 <= "111111111100110110100000000000000000";
        when "10000000010" => n11 <= "111111111001101101100000000000000000";
        when "10000000011" => n11 <= "111111110110100100100000000000000001";
        when "10000000100" => n11 <= "111111110011011011100000000000000010";
        when "10000000101" => n11 <= "111111110000010010100000000000000011";
        when "10000000110" => n11 <= "111111101101001001100000000000000101";
        when "10000000111" => n11 <= "111111101010000000100000000000000111";
        when "10000001000" => n11 <= "111111100110110111100000000000001001";
        when "10000001001" => n11 <= "111111100011101110100000000000001100";
        when "10000001010" => n11 <= "111111100000100101100000000000001111";
        when "10000001011" => n11 <= "111111011101011100100000000000010010";
        when "10000001100" => n11 <= "111111011010010011100000000000010110";
        when "10000001101" => n11 <= "111111010111001010100000000000011010";
        when "10000001110" => n11 <= "111111010100000001100000000000011110";
        when "10000001111" => n11 <= "111111010000111000100000000000100010";
        when "10000010000" => n11 <= "111111001101101111100000000000100111";
        when "10000010001" => n11 <= "111111001010100110100000000000101100";
        when "10000010010" => n11 <= "111111000111011101100000000000110001";
        when "10000010011" => n11 <= "111111000100010100100000000000110111";
        when "10000010100" => n11 <= "111111000001001011100000000000111101";
        when "10000010101" => n11 <= "111110111110000010100000000001000100";
        when "10000010110" => n11 <= "111110111010111001100000000001001010";
        when "10000010111" => n11 <= "111110110111110000100000000001010001";
        when "10000011000" => n11 <= "111110110100100111100000000001011000";
        when "10000011001" => n11 <= "111110110001011110100000000001100000";
        when "10000011010" => n11 <= "111110101110010101100000000001101000";
        when "10000011011" => n11 <= "111110101011001100100000000001110000";
        when "10000011100" => n11 <= "111110101000000011100000000001111000";
        when "10000011101" => n11 <= "111110100100111011100000000010000001";
        when "10000011110" => n11 <= "111110100001110010100000000010001010";
        when "10000011111" => n11 <= "111110011110101001100000000010010100";
        when "10000100000" => n11 <= "111110011011100000100000000010011101";
        when "10000100001" => n11 <= "111110011000010111100000000010100111";
        when "10000100010" => n11 <= "111110010101001110100000000010110010";
        when "10000100011" => n11 <= "111110010010000110100000000010111100";
        when "10000100100" => n11 <= "111110001110111101100000000011000111";
        when "10000100101" => n11 <= "111110001011110100100000000011010011";
        when "10000100110" => n11 <= "111110001000101011100000000011011110";
        when "10000100111" => n11 <= "111110000101100011100000000011101010";
        when "10000101000" => n11 <= "111110000010011010100000000011110110";
        when "10000101001" => n11 <= "111101111111010001100000000100000011";
        when "10000101010" => n11 <= "111101111100001001100000000100001111";
        when "10000101011" => n11 <= "111101111001000000100000000100011101";
        when "10000101100" => n11 <= "111101110101110111100000000100101010";
        when "10000101101" => n11 <= "111101110010101111100000000100111000";
        when "10000101110" => n11 <= "111101101111100110100000000101000110";
        when "10000101111" => n11 <= "111101101100011110100000000101010100";
        when "10000110000" => n11 <= "111101101001010101100000000101100011";
        when "10000110001" => n11 <= "111101100110001101100000000101110010";
        when "10000110010" => n11 <= "111101100011000100100000000110000001";
        when "10000110011" => n11 <= "111101011111111100100000000110010000";
        when "10000110100" => n11 <= "111101011100110011100000000110100000";
        when "10000110101" => n11 <= "111101011001101011100000000110110000";
        when "10000110110" => n11 <= "111101010110100011100000000111000001";
        when "10000110111" => n11 <= "111101010011011010100000000111010010";
        when "10000111000" => n11 <= "111101010000010010100000000111100011";
        when "10000111001" => n11 <= "111101001101001010100000000111110100";
        when "10000111010" => n11 <= "111101001010000001100000001000000110";
        when "10000111011" => n11 <= "111101000110111001100000001000011000";
        when "10000111100" => n11 <= "111101000011110001100000001000101010";
        when "10000111101" => n11 <= "111101000000101001100000001000111101";
        when "10000111110" => n11 <= "111100111101100000100000001001010000";
        when "10000111111" => n11 <= "111100111010011000100000001001100011";
        when "10001000000" => n11 <= "111100110111010000100000001001110111";
        when "10001000001" => n11 <= "111100110100001000100000001010001011";
        when "10001000010" => n11 <= "111100110001000000100000001010011111";
        when "10001000011" => n11 <= "111100101101111000100000001010110011";
        when "10001000100" => n11 <= "111100101010110000100000001011001000";
        when "10001000101" => n11 <= "111100100111101000100000001011011101";
        when "10001000110" => n11 <= "111100100100100000100000001011110010";
        when "10001000111" => n11 <= "111100100001011000100000001100001000";
        when "10001001000" => n11 <= "111100011110010000100000001100011110";
        when "10001001001" => n11 <= "111100011011001001100000001100110100";
        when "10001001010" => n11 <= "111100011000000001100000001101001011";
        when "10001001011" => n11 <= "111100010100111001100000001101100010";
        when "10001001100" => n11 <= "111100010001110001100000001101111001";
        when "10001001101" => n11 <= "111100001110101010100000001110010001";
        when "10001001110" => n11 <= "111100001011100010100000001110101001";
        when "10001001111" => n11 <= "111100001000011010100000001111000001";
        when "10001010000" => n11 <= "111100000101010011100000001111011001";
        when "10001010001" => n11 <= "111100000010001011100000001111110010";
        when "10001010010" => n11 <= "111011111111000100100000010000001011";
        when "10001010011" => n11 <= "111011111011111100100000010000100100";
        when "10001010100" => n11 <= "111011111000110101100000010000111110";
        when "10001010101" => n11 <= "111011110101101110100000010001011000";
        when "10001010110" => n11 <= "111011110010100110100000010001110010";
        when "10001010111" => n11 <= "111011101111011111100000010010001101";
        when "10001011000" => n11 <= "111011101100011000100000010010101000";
        when "10001011001" => n11 <= "111011101001010001100000010011000011";
        when "10001011010" => n11 <= "111011100110001001100000010011011111";
        when "10001011011" => n11 <= "111011100011000010100000010011111010";
        when "10001011100" => n11 <= "111011011111111011100000010100010111";
        when "10001011101" => n11 <= "111011011100110100100000010100110011";
        when "10001011110" => n11 <= "111011011001101101100000010101010000";
        when "10001011111" => n11 <= "111011010110100110100000010101101101";
        when "10001100000" => n11 <= "111011010011011111100000010110001010";
        when "10001100001" => n11 <= "111011010000011000100000010110101000";
        when "10001100010" => n11 <= "111011001101010010100000010111000110";
        when "10001100011" => n11 <= "111011001010001011100000010111100100";
        when "10001100100" => n11 <= "111011000111000100100000011000000011";
        when "10001100101" => n11 <= "111011000011111101100000011000100001";
        when "10001100110" => n11 <= "111011000000110111100000011001000001";
        when "10001100111" => n11 <= "111010111101110000100000011001100000";
        when "10001101000" => n11 <= "111010111010101010100000011010000000";
        when "10001101001" => n11 <= "111010110111100011100000011010100000";
        when "10001101010" => n11 <= "111010110100011101100000011011000000";
        when "10001101011" => n11 <= "111010110001010110100000011011100001";
        when "10001101100" => n11 <= "111010101110010000100000011100000010";
        when "10001101101" => n11 <= "111010101011001010100000011100100011";
        when "10001101110" => n11 <= "111010101000000011100000011101000101";
        when "10001101111" => n11 <= "111010100100111101100000011101100111";
        when "10001110000" => n11 <= "111010100001110111100000011110001001";
        when "10001110001" => n11 <= "111010011110110001100000011110101100";
        when "10001110010" => n11 <= "111010011011101011100000011111001111";
        when "10001110011" => n11 <= "111010011000100101100000011111110010";
        when "10001110100" => n11 <= "111010010101011111100000100000010101";
        when "10001110101" => n11 <= "111010010010011001100000100000111001";
        when "10001110110" => n11 <= "111010001111010100100000100001011101";
        when "10001110111" => n11 <= "111010001100001110100000100010000001";
        when "10001111000" => n11 <= "111010001001001000100000100010100110";
        when "10001111001" => n11 <= "111010000110000010100000100011001011";
        when "10001111010" => n11 <= "111010000010111101100000100011110000";
        when "10001111011" => n11 <= "111001111111110111100000100100010110";
        when "10001111100" => n11 <= "111001111100110010100000100100111100";
        when "10001111101" => n11 <= "111001111001101100100000100101100010";
        when "10001111110" => n11 <= "111001110110100111100000100110001000";
        when "10001111111" => n11 <= "111001110011100010100000100110101111";
        when "10010000000" => n11 <= "111001110000011101100000100111010110";
        when "10010000001" => n11 <= "111001101101010111100000100111111101";
        when "10010000010" => n11 <= "111001101010010010100000101000100101";
        when "10010000011" => n11 <= "111001100111001101100000101001001101";
        when "10010000100" => n11 <= "111001100100001000100000101001110101";
        when "10010000101" => n11 <= "111001100001000011100000101010011110";
        when "10010000110" => n11 <= "111001011101111111100000101011000111";
        when "10010000111" => n11 <= "111001011010111010100000101011110000";
        when "10010001000" => n11 <= "111001010111110101100000101100011001";
        when "10010001001" => n11 <= "111001010100110000100000101101000011";
        when "10010001010" => n11 <= "111001010001101100100000101101101101";
        when "10010001011" => n11 <= "111001001110100111100000101110011000";
        when "10010001100" => n11 <= "111001001011100011100000101111000010";
        when "10010001101" => n11 <= "111001001000011110100000101111101101";
        when "10010001110" => n11 <= "111001000101011010100000110000011001";
        when "10010001111" => n11 <= "111001000010010110100000110001000100";
        when "10010010000" => n11 <= "111000111111010001100000110001110000";
        when "10010010001" => n11 <= "111000111100001101100000110010011100";
        when "10010010010" => n11 <= "111000111001001001100000110011001001";
        when "10010010011" => n11 <= "111000110110000101100000110011110110";
        when "10010010100" => n11 <= "111000110011000001100000110100100011";
        when "10010010101" => n11 <= "111000101111111101100000110101010000";
        when "10010010110" => n11 <= "111000101100111010100000110101111110";
        when "10010010111" => n11 <= "111000101001110110100000110110101100";
        when "10010011000" => n11 <= "111000100110110010100000110111011010";
        when "10010011001" => n11 <= "111000100011101111100000111000001001";
        when "10010011010" => n11 <= "111000100000101011100000111000111000";
        when "10010011011" => n11 <= "111000011101101000100000111001100111";
        when "10010011100" => n11 <= "111000011010100100100000111010010111";
        when "10010011101" => n11 <= "111000010111100001100000111011000110";
        when "10010011110" => n11 <= "111000010100011110100000111011110110";
        when "10010011111" => n11 <= "111000010001011011100000111100100111";
        when "10010100000" => n11 <= "111000001110011000100000111101011000";
        when "10010100001" => n11 <= "111000001011010101100000111110001001";
        when "10010100010" => n11 <= "111000001000010010100000111110111010";
        when "10010100011" => n11 <= "111000000101001111100000111111101011";
        when "10010100100" => n11 <= "111000000010001100100001000000011101";
        when "10010100101" => n11 <= "110111111111001001100001000001010000";
        when "10010100110" => n11 <= "110111111100000111100001000010000010";
        when "10010100111" => n11 <= "110111111001000100100001000010110101";
        when "10010101000" => n11 <= "110111110110000010100001000011101000";
        when "10010101001" => n11 <= "110111110010111111100001000100011011";
        when "10010101010" => n11 <= "110111101111111101100001000101001111";
        when "10010101011" => n11 <= "110111101100111011100001000110000011";
        when "10010101100" => n11 <= "110111101001111001100001000110110111";
        when "10010101101" => n11 <= "110111100110110111100001000111101100";
        when "10010101110" => n11 <= "110111100011110101100001001000100001";
        when "10010101111" => n11 <= "110111100000110011100001001001010110";
        when "10010110000" => n11 <= "110111011101110001100001001010001011";
        when "10010110001" => n11 <= "110111011010101111100001001011000001";
        when "10010110010" => n11 <= "110111010111101110100001001011110111";
        when "10010110011" => n11 <= "110111010100101100100001001100101110";
        when "10010110100" => n11 <= "110111010001101010100001001101100100";
        when "10010110101" => n11 <= "110111001110101001100001001110011011";
        when "10010110110" => n11 <= "110111001011101000100001001111010011";
        when "10010110111" => n11 <= "110111001000100111100001010000001010";
        when "10010111000" => n11 <= "110111000101100101100001010001000010";
        when "10010111001" => n11 <= "110111000010100100100001010001111010";
        when "10010111010" => n11 <= "110110111111100011100001010010110011";
        when "10010111011" => n11 <= "110110111100100010100001010011101011";
        when "10010111100" => n11 <= "110110111001100010100001010100100100";
        when "10010111101" => n11 <= "110110110110100001100001010101011110";
        when "10010111110" => n11 <= "110110110011100000100001010110010111";
        when "10010111111" => n11 <= "110110110000100000100001010111010001";
        when "10011000000" => n11 <= "110110101101011111100001011000001011";
        when "10011000001" => n11 <= "110110101010011111100001011001000110";
        when "10011000010" => n11 <= "110110100111011111100001011010000001";
        when "10011000011" => n11 <= "110110100100011110100001011010111100";
        when "10011000100" => n11 <= "110110100001011110100001011011110111";
        when "10011000101" => n11 <= "110110011110011110100001011100110011";
        when "10011000110" => n11 <= "110110011011011111100001011101101111";
        when "10011000111" => n11 <= "110110011000011111100001011110101011";
        when "10011001000" => n11 <= "110110010101011111100001011111101000";
        when "10011001001" => n11 <= "110110010010011111100001100000100101";
        when "10011001010" => n11 <= "110110001111100000100001100001100010";
        when "10011001011" => n11 <= "110110001100100000100001100010011111";
        when "10011001100" => n11 <= "110110001001100001100001100011011101";
        when "10011001101" => n11 <= "110110000110100010100001100100011011";
        when "10011001110" => n11 <= "110110000011100011100001100101011001";
        when "10011001111" => n11 <= "110110000000100100100001100110011000";
        when "10011010000" => n11 <= "110101111101100101100001100111010111";
        when "10011010001" => n11 <= "110101111010100110100001101000010110";
        when "10011010010" => n11 <= "110101110111100111100001101001010110";
        when "10011010011" => n11 <= "110101110100101000100001101010010101";
        when "10011010100" => n11 <= "110101110001101010100001101011010110";
        when "10011010101" => n11 <= "110101101110101011100001101100010110";
        when "10011010110" => n11 <= "110101101011101101100001101101010111";
        when "10011010111" => n11 <= "110101101000101111100001101110011000";
        when "10011011000" => n11 <= "110101100101110000100001101111011001";
        when "10011011001" => n11 <= "110101100010110010100001110000011010";
        when "10011011010" => n11 <= "110101011111110100100001110001011100";
        when "10011011011" => n11 <= "110101011100110111100001110010011110";
        when "10011011100" => n11 <= "110101011001111001100001110011100001";
        when "10011011101" => n11 <= "110101010110111011100001110100100100";
        when "10011011110" => n11 <= "110101010011111101100001110101100111";
        when "10011011111" => n11 <= "110101010001000000100001110110101010";
        when "10011100000" => n11 <= "110101001110000011100001110111101101";
        when "10011100001" => n11 <= "110101001011000101100001111000110001";
        when "10011100010" => n11 <= "110101001000001000100001111001110101";
        when "10011100011" => n11 <= "110101000101001011100001111010111010";
        when "10011100100" => n11 <= "110101000010001110100001111011111111";
        when "10011100101" => n11 <= "110100111111010001100001111101000100";
        when "10011100110" => n11 <= "110100111100010101100001111110001001";
        when "10011100111" => n11 <= "110100111001011000100001111111001111";
        when "10011101000" => n11 <= "110100110110011100100010000000010101";
        when "10011101001" => n11 <= "110100110011011111100010000001011011";
        when "10011101010" => n11 <= "110100110000100011100010000010100001";
        when "10011101011" => n11 <= "110100101101100111100010000011101000";
        when "10011101100" => n11 <= "110100101010101011100010000100101111";
        when "10011101101" => n11 <= "110100100111101111100010000101110110";
        when "10011101110" => n11 <= "110100100100110011100010000110111110";
        when "10011101111" => n11 <= "110100100001110111100010001000000110";
        when "10011110000" => n11 <= "110100011110111011100010001001001110";
        when "10011110001" => n11 <= "110100011100000000100010001010010111";
        when "10011110010" => n11 <= "110100011001000100100010001011100000";
        when "10011110011" => n11 <= "110100010110001001100010001100101001";
        when "10011110100" => n11 <= "110100010011001110100010001101110010";
        when "10011110101" => n11 <= "110100010000010011100010001110111100";
        when "10011110110" => n11 <= "110100001101011000100010010000000110";
        when "10011110111" => n11 <= "110100001010011101100010010001010000";
        when "10011111000" => n11 <= "110100000111100010100010010010011010";
        when "10011111001" => n11 <= "110100000100101000100010010011100101";
        when "10011111010" => n11 <= "110100000001101101100010010100110000";
        when "10011111011" => n11 <= "110011111110110011100010010101111100";
        when "10011111100" => n11 <= "110011111011111000100010010111000111";
        when "10011111101" => n11 <= "110011111000111110100010011000010011";
        when "10011111110" => n11 <= "110011110110000100100010011001011111";
        when "10011111111" => n11 <= "110011110011001010100010011010101100";
        when "10100000000" => n11 <= "110011110000010000100010011011111001";
        when "10100000001" => n11 <= "110011101101010111100010011101000110";
        when "10100000010" => n11 <= "110011101010011101100010011110010011";
        when "10100000011" => n11 <= "110011100111100100100010011111100001";
        when "10100000100" => n11 <= "110011100100101010100010100000101111";
        when "10100000101" => n11 <= "110011100001110001100010100001111101";
        when "10100000110" => n11 <= "110011011110111000100010100011001100";
        when "10100000111" => n11 <= "110011011011111111100010100100011010";
        when "10100001000" => n11 <= "110011011001000110100010100101101001";
        when "10100001001" => n11 <= "110011010110001101100010100110111001";
        when "10100001010" => n11 <= "110011010011010101100010101000001000";
        when "10100001011" => n11 <= "110011010000011100100010101001011000";
        when "10100001100" => n11 <= "110011001101100100100010101010101001";
        when "10100001101" => n11 <= "110011001010101100100010101011111001";
        when "10100001110" => n11 <= "110011000111110100100010101101001010";
        when "10100001111" => n11 <= "110011000100111100100010101110011011";
        when "10100010000" => n11 <= "110011000010000100100010101111101100";
        when "10100010001" => n11 <= "110010111111001100100010110000111110";
        when "10100010010" => n11 <= "110010111100010100100010110010010000";
        when "10100010011" => n11 <= "110010111001011101100010110011100010";
        when "10100010100" => n11 <= "110010110110100101100010110100110100";
        when "10100010101" => n11 <= "110010110011101110100010110110000111";
        when "10100010110" => n11 <= "110010110000110111100010110111011010";
        when "10100010111" => n11 <= "110010101110000000100010111000101101";
        when "10100011000" => n11 <= "110010101011001001100010111010000001";
        when "10100011001" => n11 <= "110010101000010011100010111011010101";
        when "10100011010" => n11 <= "110010100101011100100010111100101001";
        when "10100011011" => n11 <= "110010100010100101100010111101111101";
        when "10100011100" => n11 <= "110010011111101111100010111111010010";
        when "10100011101" => n11 <= "110010011100111001100011000000100111";
        when "10100011110" => n11 <= "110010011010000011100011000001111100";
        when "10100011111" => n11 <= "110010010111001101100011000011010010";
        when "10100100000" => n11 <= "110010010100010111100011000100101000";
        when "10100100001" => n11 <= "110010010001100001100011000101111110";
        when "10100100010" => n11 <= "110010001110101100100011000111010100";
        when "10100100011" => n11 <= "110010001011110110100011001000101011";
        when "10100100100" => n11 <= "110010001001000001100011001010000010";
        when "10100100101" => n11 <= "110010000110001100100011001011011001";
        when "10100100110" => n11 <= "110010000011010111100011001100110001";
        when "10100100111" => n11 <= "110010000000100010100011001110001000";
        when "10100101000" => n11 <= "110001111101101101100011001111100000";
        when "10100101001" => n11 <= "110001111010111001100011010000111001";
        when "10100101010" => n11 <= "110001111000000100100011010010010001";
        when "10100101011" => n11 <= "110001110101010000100011010011101010";
        when "10100101100" => n11 <= "110001110010011100100011010101000011";
        when "10100101101" => n11 <= "110001101111100111100011010110011101";
        when "10100101110" => n11 <= "110001101100110100100011010111110111";
        when "10100101111" => n11 <= "110001101010000000100011011001010001";
        when "10100110000" => n11 <= "110001100111001100100011011010101011";
        when "10100110001" => n11 <= "110001100100011001100011011100000101";
        when "10100110010" => n11 <= "110001100001100101100011011101100000";
        when "10100110011" => n11 <= "110001011110110010100011011110111011";
        when "10100110100" => n11 <= "110001011011111111100011100000010111";
        when "10100110101" => n11 <= "110001011001001100100011100001110010";
        when "10100110110" => n11 <= "110001010110011001100011100011001110";
        when "10100110111" => n11 <= "110001010011100110100011100100101010";
        when "10100111000" => n11 <= "110001010000110100100011100110000111";
        when "10100111001" => n11 <= "110001001110000001100011100111100100";
        when "10100111010" => n11 <= "110001001011001111100011101001000001";
        when "10100111011" => n11 <= "110001001000011101100011101010011110";
        when "10100111100" => n11 <= "110001000101101011100011101011111011";
        when "10100111101" => n11 <= "110001000010111001100011101101011001";
        when "10100111110" => n11 <= "110001000000001000100011101110110111";
        when "10100111111" => n11 <= "110000111101010110100011110000010110";
        when "10101000000" => n11 <= "110000111010100101100011110001110100";
        when "10101000001" => n11 <= "110000110111110011100011110011010011";
        when "10101000010" => n11 <= "110000110101000010100011110100110010";
        when "10101000011" => n11 <= "110000110010010001100011110110010010";
        when "10101000100" => n11 <= "110000101111100000100011110111110010";
        when "10101000101" => n11 <= "110000101100110000100011111001010010";
        when "10101000110" => n11 <= "110000101001111111100011111010110010";
        when "10101000111" => n11 <= "110000100111001111100011111100010010";
        when "10101001000" => n11 <= "110000100100011111100011111101110011";
        when "10101001001" => n11 <= "110000100001101111100011111111010100";
        when "10101001010" => n11 <= "110000011110111111100100000000110110";
        when "10101001011" => n11 <= "110000011100001111100100000010010111";
        when "10101001100" => n11 <= "110000011001011111100100000011111001";
        when "10101001101" => n11 <= "110000010110110000100100000101011011";
        when "10101001110" => n11 <= "110000010100000001100100000110111110";
        when "10101001111" => n11 <= "110000010001010001100100001000100000";
        when "10101010000" => n11 <= "110000001110100010100100001010000011";
        when "10101010001" => n11 <= "110000001011110011100100001011100111";
        when "10101010010" => n11 <= "110000001001000101100100001101001010";
        when "10101010011" => n11 <= "110000000110010110100100001110101110";
        when "10101010100" => n11 <= "110000000011101000100100010000010010";
        when "10101010101" => n11 <= "110000000000111010100100010001110110";
        when "10101010110" => n11 <= "101111111110001011100100010011011011";
        when "10101010111" => n11 <= "101111111011011110100100010101000000";
        when "10101011000" => n11 <= "101111111000110000100100010110100101";
        when "10101011001" => n11 <= "101111110110000010100100011000001010";
        when "10101011010" => n11 <= "101111110011010101100100011001110000";
        when "10101011011" => n11 <= "101111110000100111100100011011010110";
        when "10101011100" => n11 <= "101111101101111010100100011100111100";
        when "10101011101" => n11 <= "101111101011001101100100011110100010";
        when "10101011110" => n11 <= "101111101000100000100100100000001001";
        when "10101011111" => n11 <= "101111100101110100100100100001110000";
        when "10101100000" => n11 <= "101111100011000111100100100011010111";
        when "10101100001" => n11 <= "101111100000011011100100100100111111";
        when "10101100010" => n11 <= "101111011101101110100100100110100111";
        when "10101100011" => n11 <= "101111011011000010100100101000001111";
        when "10101100100" => n11 <= "101111011000010110100100101001110111";
        when "10101100101" => n11 <= "101111010101101011100100101011011111";
        when "10101100110" => n11 <= "101111010010111111100100101101001000";
        when "10101100111" => n11 <= "101111010000010100100100101110110001";
        when "10101101000" => n11 <= "101111001101101000100100110000011011";
        when "10101101001" => n11 <= "101111001010111101100100110010000100";
        when "10101101010" => n11 <= "101111001000010010100100110011101110";
        when "10101101011" => n11 <= "101111000101101000100100110101011000";
        when "10101101100" => n11 <= "101111000010111101100100110111000011";
        when "10101101101" => n11 <= "101111000000010011100100111000101101";
        when "10101101110" => n11 <= "101110111101101000100100111010011000";
        when "10101101111" => n11 <= "101110111010111110100100111100000011";
        when "10101110000" => n11 <= "101110111000010100100100111101101111";
        when "10101110001" => n11 <= "101110110101101011100100111111011011";
        when "10101110010" => n11 <= "101110110011000001100101000001000111";
        when "10101110011" => n11 <= "101110110000010111100101000010110011";
        when "10101110100" => n11 <= "101110101101101110100101000100011111";
        when "10101110101" => n11 <= "101110101011000101100101000110001100";
        when "10101110110" => n11 <= "101110101000011100100101000111111001";
        when "10101110111" => n11 <= "101110100101110011100101001001100110";
        when "10101111000" => n11 <= "101110100011001011100101001011010100";
        when "10101111001" => n11 <= "101110100000100010100101001101000001";
        when "10101111010" => n11 <= "101110011101111010100101001110110000";
        when "10101111011" => n11 <= "101110011011010010100101010000011110";
        when "10101111100" => n11 <= "101110011000101010100101010010001100";
        when "10101111101" => n11 <= "101110010110000010100101010011111011";
        when "10101111110" => n11 <= "101110010011011010100101010101101010";
        when "10101111111" => n11 <= "101110010000110011100101010111011010";
        when "10110000000" => n11 <= "101110001110001100100101011001001001";
        when "10110000001" => n11 <= "101110001011100101100101011010111001";
        when "10110000010" => n11 <= "101110001000111110100101011100101001";
        when "10110000011" => n11 <= "101110000110010111100101011110011001";
        when "10110000100" => n11 <= "101110000011110000100101100000001010";
        when "10110000101" => n11 <= "101110000001001010100101100001111011";
        when "10110000110" => n11 <= "101101111110100100100101100011101100";
        when "10110000111" => n11 <= "101101111011111110100101100101011101";
        when "10110001000" => n11 <= "101101111001011000100101100111001111";
        when "10110001001" => n11 <= "101101110110110010100101101001000001";
        when "10110001010" => n11 <= "101101110100001101100101101010110011";
        when "10110001011" => n11 <= "101101110001100111100101101100100101";
        when "10110001100" => n11 <= "101101101111000010100101101110011000";
        when "10110001101" => n11 <= "101101101100011101100101110000001011";
        when "10110001110" => n11 <= "101101101001111000100101110001111110";
        when "10110001111" => n11 <= "101101100111010100100101110011110001";
        when "10110010000" => n11 <= "101101100100101111100101110101100101";
        when "10110010001" => n11 <= "101101100010001011100101110111011001";
        when "10110010010" => n11 <= "101101011111100111100101111001001101";
        when "10110010011" => n11 <= "101101011101000011100101111011000001";
        when "10110010100" => n11 <= "101101011010011111100101111100110110";
        when "10110010101" => n11 <= "101101010111111011100101111110101011";
        when "10110010110" => n11 <= "101101010101011000100110000000100000";
        when "10110010111" => n11 <= "101101010010110101100110000010010110";
        when "10110011000" => n11 <= "101101010000010010100110000100001011";
        when "10110011001" => n11 <= "101101001101101111100110000110000001";
        when "10110011010" => n11 <= "101101001011001100100110000111110111";
        when "10110011011" => n11 <= "101101001000101010100110001001101110";
        when "10110011100" => n11 <= "101101000110000111100110001011100100";
        when "10110011101" => n11 <= "101101000011100101100110001101011011";
        when "10110011110" => n11 <= "101101000001000011100110001111010010";
        when "10110011111" => n11 <= "101100111110100010100110010001001010";
        when "10110100000" => n11 <= "101100111100000000100110010011000001";
        when "10110100001" => n11 <= "101100111001011111100110010100111001";
        when "10110100010" => n11 <= "101100110110111101100110010110110010";
        when "10110100011" => n11 <= "101100110100011100100110011000101010";
        when "10110100100" => n11 <= "101100110001111011100110011010100011";
        when "10110100101" => n11 <= "101100101111011011100110011100011011";
        when "10110100110" => n11 <= "101100101100111010100110011110010101";
        when "10110100111" => n11 <= "101100101010011010100110100000001110";
        when "10110101000" => n11 <= "101100100111111010100110100010001000";
        when "10110101001" => n11 <= "101100100101011010100110100100000001";
        when "10110101010" => n11 <= "101100100010111010100110100101111100";
        when "10110101011" => n11 <= "101100100000011011100110100111110110";
        when "10110101100" => n11 <= "101100011101111011100110101001110001";
        when "10110101101" => n11 <= "101100011011011100100110101011101011";
        when "10110101110" => n11 <= "101100011000111101100110101101100110";
        when "10110101111" => n11 <= "101100010110011110100110101111100010";
        when "10110110000" => n11 <= "101100010100000000100110110001011101";
        when "10110110001" => n11 <= "101100010001100001100110110011011001";
        when "10110110010" => n11 <= "101100001111000011100110110101010101";
        when "10110110011" => n11 <= "101100001100100101100110110111010010";
        when "10110110100" => n11 <= "101100001010000111100110111001001110";
        when "10110110101" => n11 <= "101100000111101010100110111011001011";
        when "10110110110" => n11 <= "101100000101001100100110111101001000";
        when "10110110111" => n11 <= "101100000010101111100110111111000101";
        when "10110111000" => n11 <= "101100000000010010100111000001000011";
        when "10110111001" => n11 <= "101011111101110101100111000011000000";
        when "10110111010" => n11 <= "101011111011011000100111000100111110";
        when "10110111011" => n11 <= "101011111000111100100111000110111101";
        when "10110111100" => n11 <= "101011110110100000100111001000111011";
        when "10110111101" => n11 <= "101011110100000011100111001010111010";
        when "10110111110" => n11 <= "101011110001101000100111001100111001";
        when "10110111111" => n11 <= "101011101111001100100111001110111000";
        when "10111000000" => n11 <= "101011101100110000100111010000110111";
        when "10111000001" => n11 <= "101011101010010101100111010010110111";
        when "10111000010" => n11 <= "101011100111111010100111010100110111";
        when "10111000011" => n11 <= "101011100101011111100111010110110111";
        when "10111000100" => n11 <= "101011100011000100100111011000111000";
        when "10111000101" => n11 <= "101011100000101010100111011010111000";
        when "10111000110" => n11 <= "101011011110001111100111011100111001";
        when "10111000111" => n11 <= "101011011011110101100111011110111010";
        when "10111001000" => n11 <= "101011011001011011100111100000111011";
        when "10111001001" => n11 <= "101011010111000001100111100010111101";
        when "10111001010" => n11 <= "101011010100101000100111100100111111";
        when "10111001011" => n11 <= "101011010010001111100111100111000001";
        when "10111001100" => n11 <= "101011001111110101100111101001000011";
        when "10111001101" => n11 <= "101011001101011100100111101011000110";
        when "10111001110" => n11 <= "101011001011000100100111101101001000";
        when "10111001111" => n11 <= "101011001000101011100111101111001011";
        when "10111010000" => n11 <= "101011000110010011100111110001001111";
        when "10111010001" => n11 <= "101011000011111011100111110011010010";
        when "10111010010" => n11 <= "101011000001100011100111110101010110";
        when "10111010011" => n11 <= "101010111111001011100111110111011010";
        when "10111010100" => n11 <= "101010111100110011100111111001011110";
        when "10111010101" => n11 <= "101010111010011100100111111011100010";
        when "10111010110" => n11 <= "101010111000000101100111111101100111";
        when "10111010111" => n11 <= "101010110101101110100111111111101100";
        when "10111011000" => n11 <= "101010110011010111101000000001110001";
        when "10111011001" => n11 <= "101010110001000001101000000011110110";
        when "10111011010" => n11 <= "101010101110101011101000000101111100";
        when "10111011011" => n11 <= "101010101100010100101000001000000001";
        when "10111011100" => n11 <= "101010101001111110101000001010000111";
        when "10111011101" => n11 <= "101010100111101001101000001100001110";
        when "10111011110" => n11 <= "101010100101010011101000001110010100";
        when "10111011111" => n11 <= "101010100010111110101000010000011011";
        when "10111100000" => n11 <= "101010100000101001101000010010100010";
        when "10111100001" => n11 <= "101010011110010100101000010100101001";
        when "10111100010" => n11 <= "101010011011111111101000010110110000";
        when "10111100011" => n11 <= "101010011001101011101000011000111000";
        when "10111100100" => n11 <= "101010010111010111101000011010111111";
        when "10111100101" => n11 <= "101010010101000011101000011101001000";
        when "10111100110" => n11 <= "101010010010101111101000011111010000";
        when "10111100111" => n11 <= "101010010000011011101000100001011000";
        when "10111101000" => n11 <= "101010001110001000101000100011100001";
        when "10111101001" => n11 <= "101010001011110101101000100101101010";
        when "10111101010" => n11 <= "101010001001100010101000100111110011";
        when "10111101011" => n11 <= "101010000111001111101000101001111101";
        when "10111101100" => n11 <= "101010000100111100101000101100000110";
        when "10111101101" => n11 <= "101010000010101010101000101110010000";
        when "10111101110" => n11 <= "101010000000011000101000110000011010";
        when "10111101111" => n11 <= "101001111110000110101000110010100100";
        when "10111110000" => n11 <= "101001111011110100101000110100101111";
        when "10111110001" => n11 <= "101001111001100011101000110110111010";
        when "10111110010" => n11 <= "101001110111010001101000111001000101";
        when "10111110011" => n11 <= "101001110101000000101000111011010000";
        when "10111110100" => n11 <= "101001110010101111101000111101011011";
        when "10111110101" => n11 <= "101001110000011111101000111111100111";
        when "10111110110" => n11 <= "101001101110001110101001000001110011";
        when "10111110111" => n11 <= "101001101011111110101001000011111111";
        when "10111111000" => n11 <= "101001101001101110101001000110001011";
        when "10111111001" => n11 <= "101001100111011110101001001000011000";
        when "10111111010" => n11 <= "101001100101001111101001001010100101";
        when "10111111011" => n11 <= "101001100010111111101001001100110001";
        when "10111111100" => n11 <= "101001100000110000101001001110111111";
        when "10111111101" => n11 <= "101001011110100001101001010001001100";
        when "10111111110" => n11 <= "101001011100010010101001010011011010";
        when "10111111111" => n11 <= "101001011010000100101001010101101000";
        when "11000000000" => n11 <= "101001010111110110101001010111110110";
        when "11000000001" => n11 <= "101001010101101000101001011010000100";
        when "11000000010" => n11 <= "101001010011011010101001011100010010";
        when "11000000011" => n11 <= "101001010001001100101001011110100001";
        when "11000000100" => n11 <= "101001001110111111101001100000110000";
        when "11000000101" => n11 <= "101001001100110001101001100010111111";
        when "11000000110" => n11 <= "101001001010100101101001100101001111";
        when "11000000111" => n11 <= "101001001000011000101001100111011110";
        when "11000001000" => n11 <= "101001000110001011101001101001101110";
        when "11000001001" => n11 <= "101001000011111111101001101011111110";
        when "11000001010" => n11 <= "101001000001110011101001101110001110";
        when "11000001011" => n11 <= "101000111111100111101001110000011111";
        when "11000001100" => n11 <= "101000111101011011101001110010101111";
        when "11000001101" => n11 <= "101000111011010000101001110101000000";
        when "11000001110" => n11 <= "101000111001000101101001110111010001";
        when "11000001111" => n11 <= "101000110110111010101001111001100011";
        when "11000010000" => n11 <= "101000110100101111101001111011110100";
        when "11000010001" => n11 <= "101000110010100100101001111110000110";
        when "11000010010" => n11 <= "101000110000011010101010000000011000";
        when "11000010011" => n11 <= "101000101110010000101010000010101010";
        when "11000010100" => n11 <= "101000101100000110101010000100111100";
        when "11000010101" => n11 <= "101000101001111101101010000111001111";
        when "11000010110" => n11 <= "101000100111110011101010001001100010";
        when "11000010111" => n11 <= "101000100101101010101010001011110101";
        when "11000011000" => n11 <= "101000100011100001101010001110001000";
        when "11000011001" => n11 <= "101000100001011000101010010000011011";
        when "11000011010" => n11 <= "101000011111010000101010010010101111";
        when "11000011011" => n11 <= "101000011101001000101010010101000011";
        when "11000011100" => n11 <= "101000011010111111101010010111010111";
        when "11000011101" => n11 <= "101000011000111000101010011001101011";
        when "11000011110" => n11 <= "101000010110110000101010011011111111";
        when "11000011111" => n11 <= "101000010100101001101010011110010100";
        when "11000100000" => n11 <= "101000010010100010101010100000101001";
        when "11000100001" => n11 <= "101000010000011011101010100010111110";
        when "11000100010" => n11 <= "101000001110010100101010100101010011";
        when "11000100011" => n11 <= "101000001100001110101010100111101001";
        when "11000100100" => n11 <= "101000001010000111101010101001111110";
        when "11000100101" => n11 <= "101000001000000001101010101100010100";
        when "11000100110" => n11 <= "101000000101111100101010101110101011";
        when "11000100111" => n11 <= "101000000011110110101010110001000001";
        when "11000101000" => n11 <= "101000000001110001101010110011010111";
        when "11000101001" => n11 <= "100111111111101100101010110101101110";
        when "11000101010" => n11 <= "100111111101100111101010111000000101";
        when "11000101011" => n11 <= "100111111011100010101010111010011100";
        when "11000101100" => n11 <= "100111111001011110101010111100110011";
        when "11000101101" => n11 <= "100111110111011010101010111111001011";
        when "11000101110" => n11 <= "100111110101010110101011000001100011";
        when "11000101111" => n11 <= "100111110011010010101011000011111011";
        when "11000110000" => n11 <= "100111110001001111101011000110010011";
        when "11000110001" => n11 <= "100111101111001011101011001000101011";
        when "11000110010" => n11 <= "100111101101001000101011001011000100";
        when "11000110011" => n11 <= "100111101011000110101011001101011100";
        when "11000110100" => n11 <= "100111101001000011101011001111110101";
        when "11000110101" => n11 <= "100111100111000001101011010010001111";
        when "11000110110" => n11 <= "100111100100111111101011010100101000";
        when "11000110111" => n11 <= "100111100010111101101011010111000001";
        when "11000111000" => n11 <= "100111100000111011101011011001011011";
        when "11000111001" => n11 <= "100111011110111010101011011011110101";
        when "11000111010" => n11 <= "100111011100111001101011011110001111";
        when "11000111011" => n11 <= "100111011010111000101011100000101010";
        when "11000111100" => n11 <= "100111011000111000101011100011000100";
        when "11000111101" => n11 <= "100111010110110111101011100101011111";
        when "11000111110" => n11 <= "100111010100110111101011100111111010";
        when "11000111111" => n11 <= "100111010010110111101011101010010101";
        when "11001000000" => n11 <= "100111010000110111101011101100110000";
        when "11001000001" => n11 <= "100111001110111000101011101111001100";
        when "11001000010" => n11 <= "100111001100111001101011110001101000";
        when "11001000011" => n11 <= "100111001010111010101011110100000011";
        when "11001000100" => n11 <= "100111001000111011101011110110100000";
        when "11001000101" => n11 <= "100111000110111101101011111000111100";
        when "11001000110" => n11 <= "100111000100111110101011111011011000";
        when "11001000111" => n11 <= "100111000011000000101011111101110101";
        when "11001001000" => n11 <= "100111000001000011101100000000010010";
        when "11001001001" => n11 <= "100110111111000101101100000010101111";
        when "11001001010" => n11 <= "100110111101001000101100000101001100";
        when "11001001011" => n11 <= "100110111011001011101100000111101010";
        when "11001001100" => n11 <= "100110111001001110101100001010000111";
        when "11001001101" => n11 <= "100110110111010010101100001100100101";
        when "11001001110" => n11 <= "100110110101010101101100001111000011";
        when "11001001111" => n11 <= "100110110011011001101100010001100001";
        when "11001010000" => n11 <= "100110110001011101101100010100000000";
        when "11001010001" => n11 <= "100110101111100010101100010110011110";
        when "11001010010" => n11 <= "100110101101100110101100011000111101";
        when "11001010011" => n11 <= "100110101011101011101100011011011100";
        when "11001010100" => n11 <= "100110101001110001101100011101111011";
        when "11001010101" => n11 <= "100110100111110110101100100000011011";
        when "11001010110" => n11 <= "100110100101111100101100100010111010";
        when "11001010111" => n11 <= "100110100100000001101100100101011010";
        when "11001011000" => n11 <= "100110100010001000101100100111111010";
        when "11001011001" => n11 <= "100110100000001110101100101010011010";
        when "11001011010" => n11 <= "100110011110010101101100101100111010";
        when "11001011011" => n11 <= "100110011100011011101100101111011011";
        when "11001011100" => n11 <= "100110011010100011101100110001111011";
        when "11001011101" => n11 <= "100110011000101010101100110100011100";
        when "11001011110" => n11 <= "100110010110110010101100110110111101";
        when "11001011111" => n11 <= "100110010100111001101100111001011111";
        when "11001100000" => n11 <= "100110010011000001101100111100000000";
        when "11001100001" => n11 <= "100110010001001010101100111110100010";
        when "11001100010" => n11 <= "100110001111010010101101000001000011";
        when "11001100011" => n11 <= "100110001101011011101101000011100101";
        when "11001100100" => n11 <= "100110001011100100101101000110000111";
        when "11001100101" => n11 <= "100110001001101110101101001000101010";
        when "11001100110" => n11 <= "100110000111110111101101001011001100";
        when "11001100111" => n11 <= "100110000110000001101101001101101111";
        when "11001101000" => n11 <= "100110000100001011101101010000010010";
        when "11001101001" => n11 <= "100110000010010110101101010010110101";
        when "11001101010" => n11 <= "100110000000100000101101010101011000";
        when "11001101011" => n11 <= "100101111110101011101101010111111011";
        when "11001101100" => n11 <= "100101111100110110101101011010011111";
        when "11001101101" => n11 <= "100101111011000001101101011101000011";
        when "11001101110" => n11 <= "100101111001001101101101011111100111";
        when "11001101111" => n11 <= "100101110111011001101101100010001011";
        when "11001110000" => n11 <= "100101110101100101101101100100101111";
        when "11001110001" => n11 <= "100101110011110001101101100111010100";
        when "11001110010" => n11 <= "100101110001111110101101101001111000";
        when "11001110011" => n11 <= "100101110000001011101101101100011101";
        when "11001110100" => n11 <= "100101101110011000101101101111000010";
        when "11001110101" => n11 <= "100101101100100101101101110001100111";
        when "11001110110" => n11 <= "100101101010110011101101110100001101";
        when "11001110111" => n11 <= "100101101001000001101101110110110010";
        when "11001111000" => n11 <= "100101100111001111101101111001011000";
        when "11001111001" => n11 <= "100101100101011101101101111011111110";
        when "11001111010" => n11 <= "100101100011101100101101111110100100";
        when "11001111011" => n11 <= "100101100001111011101110000001001010";
        when "11001111100" => n11 <= "100101100000001010101110000011110000";
        when "11001111101" => n11 <= "100101011110011001101110000110010111";
        when "11001111110" => n11 <= "100101011100101001101110001000111110";
        when "11001111111" => n11 <= "100101011010111001101110001011100101";
        when "11010000000" => n11 <= "100101011001001001101110001110001100";
        when "11010000001" => n11 <= "100101010111011010101110010000110011";
        when "11010000010" => n11 <= "100101010101101010101110010011011010";
        when "11010000011" => n11 <= "100101010011111011101110010110000010";
        when "11010000100" => n11 <= "100101010010001100101110011000101010";
        when "11010000101" => n11 <= "100101010000011110101110011011010010";
        when "11010000110" => n11 <= "100101001110110000101110011101111010";
        when "11010000111" => n11 <= "100101001101000001101110100000100010";
        when "11010001000" => n11 <= "100101001011010100101110100011001011";
        when "11010001001" => n11 <= "100101001001100110101110100101110011";
        when "11010001010" => n11 <= "100101000111111001101110101000011100";
        when "11010001011" => n11 <= "100101000110001100101110101011000101";
        when "11010001100" => n11 <= "100101000100011111101110101101101110";
        when "11010001101" => n11 <= "100101000010110011101110110000010111";
        when "11010001110" => n11 <= "100101000001000111101110110011000001";
        when "11010001111" => n11 <= "100100111111011011101110110101101011";
        when "11010010000" => n11 <= "100100111101101111101110111000010100";
        when "11010010001" => n11 <= "100100111100000011101110111010111110";
        when "11010010010" => n11 <= "100100111010011000101110111101101000";
        when "11010010011" => n11 <= "100100111000101101101111000000010011";
        when "11010010100" => n11 <= "100100110111000011101111000010111101";
        when "11010010101" => n11 <= "100100110101011000101111000101101000";
        when "11010010110" => n11 <= "100100110011101110101111001000010010";
        when "11010010111" => n11 <= "100100110010000100101111001010111101";
        when "11010011000" => n11 <= "100100110000011011101111001101101000";
        when "11010011001" => n11 <= "100100101110110001101111010000010100";
        when "11010011010" => n11 <= "100100101101001000101111010010111111";
        when "11010011011" => n11 <= "100100101011011111101111010101101011";
        when "11010011100" => n11 <= "100100101001110111101111011000010110";
        when "11010011101" => n11 <= "100100101000001111101111011011000010";
        when "11010011110" => n11 <= "100100100110100111101111011101101110";
        when "11010011111" => n11 <= "100100100100111111101111100000011011";
        when "11010100000" => n11 <= "100100100011010111101111100011000111";
        when "11010100001" => n11 <= "100100100001110000101111100101110100";
        when "11010100010" => n11 <= "100100100000001001101111101000100000";
        when "11010100011" => n11 <= "100100011110100010101111101011001101";
        when "11010100100" => n11 <= "100100011100111100101111101101111010";
        when "11010100101" => n11 <= "100100011011010110101111110000100111";
        when "11010100110" => n11 <= "100100011001110000101111110011010101";
        when "11010100111" => n11 <= "100100011000001010101111110110000010";
        when "11010101000" => n11 <= "100100010110100101101111111000110000";
        when "11010101001" => n11 <= "100100010101000000101111111011011110";
        when "11010101010" => n11 <= "100100010011011011101111111110001011";
        when "11010101011" => n11 <= "100100010001110110110000000000111010";
        when "11010101100" => n11 <= "100100010000010010110000000011101000";
        when "11010101101" => n11 <= "100100001110101110110000000110010110";
        when "11010101110" => n11 <= "100100001101001010110000001001000101";
        when "11010101111" => n11 <= "100100001011100111110000001011110011";
        when "11010110000" => n11 <= "100100001010000011110000001110100010";
        when "11010110001" => n11 <= "100100001000100000110000010001010001";
        when "11010110010" => n11 <= "100100000110111110110000010100000001";
        when "11010110011" => n11 <= "100100000101011011110000010110110000";
        when "11010110100" => n11 <= "100100000011111001110000011001011111";
        when "11010110101" => n11 <= "100100000010010111110000011100001111";
        when "11010110110" => n11 <= "100100000000110110110000011110111111";
        when "11010110111" => n11 <= "100011111111010100110000100001101111";
        when "11010111000" => n11 <= "100011111101110011110000100100011111";
        when "11010111001" => n11 <= "100011111100010010110000100111001111";
        when "11010111010" => n11 <= "100011111010110010110000101001111111";
        when "11010111011" => n11 <= "100011111001010010110000101100110000";
        when "11010111100" => n11 <= "100011110111110010110000101111100000";
        when "11010111101" => n11 <= "100011110110010010110000110010010001";
        when "11010111110" => n11 <= "100011110100110010110000110101000010";
        when "11010111111" => n11 <= "100011110011010011110000110111110011";
        when "11011000000" => n11 <= "100011110001110100110000111010100101";
        when "11011000001" => n11 <= "100011110000010110110000111101010110";
        when "11011000010" => n11 <= "100011101110110111110001000000001000";
        when "11011000011" => n11 <= "100011101101011001110001000010111001";
        when "11011000100" => n11 <= "100011101011111011110001000101101011";
        when "11011000101" => n11 <= "100011101010011110110001001000011101";
        when "11011000110" => n11 <= "100011101001000001110001001011001111";
        when "11011000111" => n11 <= "100011100111100100110001001110000001";
        when "11011001000" => n11 <= "100011100110000111110001010000110100";
        when "11011001001" => n11 <= "100011100100101010110001010011100110";
        when "11011001010" => n11 <= "100011100011001110110001010110011001";
        when "11011001011" => n11 <= "100011100001110010110001011001001100";
        when "11011001100" => n11 <= "100011100000010111110001011011111111";
        when "11011001101" => n11 <= "100011011110111011110001011110110010";
        when "11011001110" => n11 <= "100011011101100000110001100001100101";
        when "11011001111" => n11 <= "100011011100000101110001100100011001";
        when "11011010000" => n11 <= "100011011010101011110001100111001100";
        when "11011010001" => n11 <= "100011011001010001110001101010000000";
        when "11011010010" => n11 <= "100011010111110111110001101100110100";
        when "11011010011" => n11 <= "100011010110011101110001101111100111";
        when "11011010100" => n11 <= "100011010101000011110001110010011100";
        when "11011010101" => n11 <= "100011010011101010110001110101010000";
        when "11011010110" => n11 <= "100011010010010001110001111000000100";
        when "11011010111" => n11 <= "100011010000111001110001111010111001";
        when "11011011000" => n11 <= "100011001111100000110001111101101101";
        when "11011011001" => n11 <= "100011001110001000110010000000100010";
        when "11011011010" => n11 <= "100011001100110001110010000011010111";
        when "11011011011" => n11 <= "100011001011011001110010000110001100";
        when "11011011100" => n11 <= "100011001010000010110010001001000001";
        when "11011011101" => n11 <= "100011001000101011110010001011110110";
        when "11011011110" => n11 <= "100011000111010100110010001110101100";
        when "11011011111" => n11 <= "100011000101111110110010010001100001";
        when "11011100000" => n11 <= "100011000100101000110010010100010111";
        when "11011100001" => n11 <= "100011000011010010110010010111001101";
        when "11011100010" => n11 <= "100011000001111100110010011010000011";
        when "11011100011" => n11 <= "100011000000100111110010011100111001";
        when "11011100100" => n11 <= "100010111111010010110010011111101111";
        when "11011100101" => n11 <= "100010111101111101110010100010100101";
        when "11011100110" => n11 <= "100010111100101001110010100101011100";
        when "11011100111" => n11 <= "100010111011010101110010101000010011";
        when "11011101000" => n11 <= "100010111010000001110010101011001001";
        when "11011101001" => n11 <= "100010111000101101110010101110000000";
        when "11011101010" => n11 <= "100010110111011010110010110000110111";
        when "11011101011" => n11 <= "100010110110000111110010110011101110";
        when "11011101100" => n11 <= "100010110100110100110010110110100101";
        when "11011101101" => n11 <= "100010110011100010110010111001011101";
        when "11011101110" => n11 <= "100010110010010000110010111100010100";
        when "11011101111" => n11 <= "100010110000111110110010111111001100";
        when "11011110000" => n11 <= "100010101111101100110011000010000100";
        when "11011110001" => n11 <= "100010101110011011110011000100111100";
        when "11011110010" => n11 <= "100010101101001010110011000111110100";
        when "11011110011" => n11 <= "100010101011111001110011001010101100";
        when "11011110100" => n11 <= "100010101010101001110011001101100100";
        when "11011110101" => n11 <= "100010101001011000110011010000011100";
        when "11011110110" => n11 <= "100010101000001000110011010011010101";
        when "11011110111" => n11 <= "100010100110111001110011010110001101";
        when "11011111000" => n11 <= "100010100101101001110011011001000110";
        when "11011111001" => n11 <= "100010100100011010110011011011111111";
        when "11011111010" => n11 <= "100010100011001100110011011110111000";
        when "11011111011" => n11 <= "100010100001111101110011100001110001";
        when "11011111100" => n11 <= "100010100000101111110011100100101010";
        when "11011111101" => n11 <= "100010011111100001110011100111100100";
        when "11011111110" => n11 <= "100010011110010011110011101010011101";
        when "11011111111" => n11 <= "100010011101000110110011101101010111";
        when "11100000000" => n11 <= "100010011011111001110011110000010000";
        when "11100000001" => n11 <= "100010011010101100110011110011001010";
        when "11100000010" => n11 <= "100010011001011111110011110110000100";
        when "11100000011" => n11 <= "100010011000010011110011111000111110";
        when "11100000100" => n11 <= "100010010111000111110011111011111000";
        when "11100000101" => n11 <= "100010010101111100110011111110110011";
        when "11100000110" => n11 <= "100010010100110000110100000001101101";
        when "11100000111" => n11 <= "100010010011100101110100000100101000";
        when "11100001000" => n11 <= "100010010010011010110100000111100010";
        when "11100001001" => n11 <= "100010010001010000110100001010011101";
        when "11100001010" => n11 <= "100010010000000110110100001101011000";
        when "11100001011" => n11 <= "100010001110111100110100010000010011";
        when "11100001100" => n11 <= "100010001101110010110100010011001110";
        when "11100001101" => n11 <= "100010001100101001110100010110001001";
        when "11100001110" => n11 <= "100010001011100000110100011001000100";
        when "11100001111" => n11 <= "100010001010010111110100011100000000";
        when "11100010000" => n11 <= "100010001001001110110100011110111011";
        when "11100010001" => n11 <= "100010001000000110110100100001110111";
        when "11100010010" => n11 <= "100010000110111110110100100100110011";
        when "11100010011" => n11 <= "100010000101110110110100100111101111";
        when "11100010100" => n11 <= "100010000100101111110100101010101011";
        when "11100010101" => n11 <= "100010000011101000110100101101100111";
        when "11100010110" => n11 <= "100010000010100001110100110000100011";
        when "11100010111" => n11 <= "100010000001011011110100110011011111";
        when "11100011000" => n11 <= "100010000000010101110100110110011100";
        when "11100011001" => n11 <= "100001111111001111110100111001011000";
        when "11100011010" => n11 <= "100001111110001001110100111100010101";
        when "11100011011" => n11 <= "100001111101000100110100111111010001";
        when "11100011100" => n11 <= "100001111011111111110101000010001110";
        when "11100011101" => n11 <= "100001111010111010110101000101001011";
        when "11100011110" => n11 <= "100001111001110101110101001000001000";
        when "11100011111" => n11 <= "100001111000110001110101001011000101";
        when "11100100000" => n11 <= "100001110111101101110101001110000011";
        when "11100100001" => n11 <= "100001110110101010110101010001000000";
        when "11100100010" => n11 <= "100001110101100111110101010011111101";
        when "11100100011" => n11 <= "100001110100100100110101010110111011";
        when "11100100100" => n11 <= "100001110011100001110101011001111001";
        when "11100100101" => n11 <= "100001110010011110110101011100110111";
        when "11100100110" => n11 <= "100001110001011100110101011111110100";
        when "11100100111" => n11 <= "100001110000011010110101100010110010";
        when "11100101000" => n11 <= "100001101111011001110101100101110000";
        when "11100101001" => n11 <= "100001101110011000110101101000101111";
        when "11100101010" => n11 <= "100001101101010111110101101011101101";
        when "11100101011" => n11 <= "100001101100010110110101101110101011";
        when "11100101100" => n11 <= "100001101011010110110101110001101010";
        when "11100101101" => n11 <= "100001101010010101110101110100101000";
        when "11100101110" => n11 <= "100001101001010110110101110111100111";
        when "11100101111" => n11 <= "100001101000010110110101111010100110";
        when "11100110000" => n11 <= "100001100111010111110101111101100101";
        when "11100110001" => n11 <= "100001100110011000110110000000100100";
        when "11100110010" => n11 <= "100001100101011001110110000011100011";
        when "11100110011" => n11 <= "100001100100011011110110000110100010";
        when "11100110100" => n11 <= "100001100011011101110110001001100001";
        when "11100110101" => n11 <= "100001100010011111110110001100100000";
        when "11100110110" => n11 <= "100001100001100010110110001111100000";
        when "11100110111" => n11 <= "100001100000100101110110010010011111";
        when "11100111000" => n11 <= "100001011111101000110110010101011111";
        when "11100111001" => n11 <= "100001011110101011110110011000011111";
        when "11100111010" => n11 <= "100001011101101111110110011011011111";
        when "11100111011" => n11 <= "100001011100110011110110011110011110";
        when "11100111100" => n11 <= "100001011011110111110110100001011110";
        when "11100111101" => n11 <= "100001011010111100110110100100011110";
        when "11100111110" => n11 <= "100001011010000001110110100111011111";
        when "11100111111" => n11 <= "100001011001000110110110101010011111";
        when "11101000000" => n11 <= "100001011000001011110110101101011111";
        when "11101000001" => n11 <= "100001010111010001110110110000100000";
        when "11101000010" => n11 <= "100001010110010111110110110011100000";
        when "11101000011" => n11 <= "100001010101011110110110110110100001";
        when "11101000100" => n11 <= "100001010100100100110110111001100010";
        when "11101000101" => n11 <= "100001010011101011110110111100100010";
        when "11101000110" => n11 <= "100001010010110011110110111111100011";
        when "11101000111" => n11 <= "100001010001111010110111000010100100";
        when "11101001000" => n11 <= "100001010001000010110111000101100101";
        when "11101001001" => n11 <= "100001010000001010110111001000100111";
        when "11101001010" => n11 <= "100001001111010011110111001011101000";
        when "11101001011" => n11 <= "100001001110011011110111001110101001";
        when "11101001100" => n11 <= "100001001101100100110111010001101010";
        when "11101001101" => n11 <= "100001001100101110110111010100101100";
        when "11101001110" => n11 <= "100001001011110111110111010111101110";
        when "11101001111" => n11 <= "100001001011000001110111011010101111";
        when "11101010000" => n11 <= "100001001010001011110111011101110001";
        when "11101010001" => n11 <= "100001001001010110110111100000110011";
        when "11101010010" => n11 <= "100001001000100001110111100011110101";
        when "11101010011" => n11 <= "100001000111101100110111100110110111";
        when "11101010100" => n11 <= "100001000110110111110111101001111001";
        when "11101010101" => n11 <= "100001000110000011110111101100111011";
        when "11101010110" => n11 <= "100001000101001111110111101111111101";
        when "11101010111" => n11 <= "100001000100011011110111110010111111";
        when "11101011000" => n11 <= "100001000011101000110111110110000010";
        when "11101011001" => n11 <= "100001000010110101110111111001000100";
        when "11101011010" => n11 <= "100001000010000010110111111100000111";
        when "11101011011" => n11 <= "100001000001010000110111111111001001";
        when "11101011100" => n11 <= "100001000000011101111000000010001100";
        when "11101011101" => n11 <= "100000111111101011111000000101001111";
        when "11101011110" => n11 <= "100000111110111010111000001000010010";
        when "11101011111" => n11 <= "100000111110001001111000001011010101";
        when "11101100000" => n11 <= "100000111101011000111000001110011000";
        when "11101100001" => n11 <= "100000111100100111111000010001011011";
        when "11101100010" => n11 <= "100000111011110110111000010100011110";
        when "11101100011" => n11 <= "100000111011000110111000010111100001";
        when "11101100100" => n11 <= "100000111010010111111000011010100100";
        when "11101100101" => n11 <= "100000111001100111111000011101101000";
        when "11101100110" => n11 <= "100000111000111000111000100000101011";
        when "11101100111" => n11 <= "100000111000001001111000100011101111";
        when "11101101000" => n11 <= "100000110111011010111000100110110010";
        when "11101101001" => n11 <= "100000110110101100111000101001110110";
        when "11101101010" => n11 <= "100000110101111110111000101100111010";
        when "11101101011" => n11 <= "100000110101010000111000101111111101";
        when "11101101100" => n11 <= "100000110100100011111000110011000001";
        when "11101101101" => n11 <= "100000110011110110111000110110000101";
        when "11101101110" => n11 <= "100000110011001001111000111001001001";
        when "11101101111" => n11 <= "100000110010011100111000111100001101";
        when "11101110000" => n11 <= "100000110001110000111000111111010001";
        when "11101110001" => n11 <= "100000110001000100111001000010010110";
        when "11101110010" => n11 <= "100000110000011001111001000101011010";
        when "11101110011" => n11 <= "100000101111101101111001001000011110";
        when "11101110100" => n11 <= "100000101111000010111001001011100011";
        when "11101110101" => n11 <= "100000101110011000111001001110100111";
        when "11101110110" => n11 <= "100000101101101101111001010001101100";
        when "11101110111" => n11 <= "100000101101000011111001010100110000";
        when "11101111000" => n11 <= "100000101100011001111001010111110101";
        when "11101111001" => n11 <= "100000101011110000111001011010111010";
        when "11101111010" => n11 <= "100000101011000111111001011101111111";
        when "11101111011" => n11 <= "100000101010011110111001100001000011";
        when "11101111100" => n11 <= "100000101001110101111001100100001000";
        when "11101111101" => n11 <= "100000101001001101111001100111001101";
        when "11101111110" => n11 <= "100000101000100101111001101010010010";
        when "11101111111" => n11 <= "100000100111111101111001101101010111";
        when "11110000000" => n11 <= "100000100111010110111001110000011101";
        when "11110000001" => n11 <= "100000100110101111111001110011100010";
        when "11110000010" => n11 <= "100000100110001000111001110110100111";
        when "11110000011" => n11 <= "100000100101100010111001111001101100";
        when "11110000100" => n11 <= "100000100100111100111001111100110010";
        when "11110000101" => n11 <= "100000100100010110111001111111110111";
        when "11110000110" => n11 <= "100000100011110000111010000010111101";
        when "11110000111" => n11 <= "100000100011001011111010000110000010";
        when "11110001000" => n11 <= "100000100010100110111010001001001000";
        when "11110001001" => n11 <= "100000100010000001111010001100001110";
        when "11110001010" => n11 <= "100000100001011101111010001111010100";
        when "11110001011" => n11 <= "100000100000111001111010010010011001";
        when "11110001100" => n11 <= "100000100000010101111010010101011111";
        when "11110001101" => n11 <= "100000011111110010111010011000100101";
        when "11110001110" => n11 <= "100000011111001111111010011011101011";
        when "11110001111" => n11 <= "100000011110101100111010011110110001";
        when "11110010000" => n11 <= "100000011110001001111010100001110111";
        when "11110010001" => n11 <= "100000011101100111111010100100111101";
        when "11110010010" => n11 <= "100000011101000101111010101000000011";
        when "11110010011" => n11 <= "100000011100100011111010101011001010";
        when "11110010100" => n11 <= "100000011100000010111010101110010000";
        when "11110010101" => n11 <= "100000011011100001111010110001010110";
        when "11110010110" => n11 <= "100000011011000000111010110100011101";
        when "11110010111" => n11 <= "100000011010100000111010110111100011";
        when "11110011000" => n11 <= "100000011010000000111010111010101010";
        when "11110011001" => n11 <= "100000011001100000111010111101110000";
        when "11110011010" => n11 <= "100000011001000001111011000000110111";
        when "11110011011" => n11 <= "100000011000100001111011000011111101";
        when "11110011100" => n11 <= "100000011000000011111011000111000100";
        when "11110011101" => n11 <= "100000010111100100111011001010001011";
        when "11110011110" => n11 <= "100000010111000110111011001101010010";
        when "11110011111" => n11 <= "100000010110101000111011010000011000";
        when "11110100000" => n11 <= "100000010110001010111011010011011111";
        when "11110100001" => n11 <= "100000010101101101111011010110100110";
        when "11110100010" => n11 <= "100000010101010000111011011001101101";
        when "11110100011" => n11 <= "100000010100110011111011011100110100";
        when "11110100100" => n11 <= "100000010100010111111011011111111011";
        when "11110100101" => n11 <= "100000010011111010111011100011000010";
        when "11110100110" => n11 <= "100000010011011111111011100110001001";
        when "11110100111" => n11 <= "100000010011000011111011101001010001";
        when "11110101000" => n11 <= "100000010010101000111011101100011000";
        when "11110101001" => n11 <= "100000010010001101111011101111011111";
        when "11110101010" => n11 <= "100000010001110010111011110010100110";
        when "11110101011" => n11 <= "100000010001011000111011110101101110";
        when "11110101100" => n11 <= "100000010000111110111011111000110101";
        when "11110101101" => n11 <= "100000010000100100111011111011111100";
        when "11110101110" => n11 <= "100000010000001011111011111111000100";
        when "11110101111" => n11 <= "100000001111110010111100000010001011";
        when "11110110000" => n11 <= "100000001111011001111100000101010011";
        when "11110110001" => n11 <= "100000001111000001111100001000011010";
        when "11110110010" => n11 <= "100000001110101001111100001011100010";
        when "11110110011" => n11 <= "100000001110010001111100001110101010";
        when "11110110100" => n11 <= "100000001101111001111100010001110001";
        when "11110110101" => n11 <= "100000001101100010111100010100111001";
        when "11110110110" => n11 <= "100000001101001011111100011000000001";
        when "11110110111" => n11 <= "100000001100110100111100011011001001";
        when "11110111000" => n11 <= "100000001100011110111100011110010000";
        when "11110111001" => n11 <= "100000001100001000111100100001011000";
        when "11110111010" => n11 <= "100000001011110010111100100100100000";
        when "11110111011" => n11 <= "100000001011011101111100100111101000";
        when "11110111100" => n11 <= "100000001011001000111100101010110000";
        when "11110111101" => n11 <= "100000001010110011111100101101111000";
        when "11110111110" => n11 <= "100000001010011111111100110001000000";
        when "11110111111" => n11 <= "100000001010001011111100110100001000";
        when "11111000000" => n11 <= "100000001001110111111100110111010000";
        when "11111000001" => n11 <= "100000001001100011111100111010011000";
        when "11111000010" => n11 <= "100000001001010000111100111101100000";
        when "11111000011" => n11 <= "100000001000111101111101000000101001";
        when "11111000100" => n11 <= "100000001000101010111101000011110001";
        when "11111000101" => n11 <= "100000001000011000111101000110111001";
        when "11111000110" => n11 <= "100000001000000110111101001010000001";
        when "11111000111" => n11 <= "100000000111110100111101001101001010";
        when "11111001000" => n11 <= "100000000111100011111101010000010010";
        when "11111001001" => n11 <= "100000000111010010111101010011011010";
        when "11111001010" => n11 <= "100000000111000001111101010110100011";
        when "11111001011" => n11 <= "100000000110110000111101011001101011";
        when "11111001100" => n11 <= "100000000110100000111101011100110011";
        when "11111001101" => n11 <= "100000000110010000111101011111111100";
        when "11111001110" => n11 <= "100000000110000001111101100011000100";
        when "11111001111" => n11 <= "100000000101110010111101100110001101";
        when "11111010000" => n11 <= "100000000101100011111101101001010101";
        when "11111010001" => n11 <= "100000000101010100111101101100011110";
        when "11111010010" => n11 <= "100000000101000110111101101111100110";
        when "11111010011" => n11 <= "100000000100111000111101110010101111";
        when "11111010100" => n11 <= "100000000100101010111101110101110111";
        when "11111010101" => n11 <= "100000000100011101111101111001000000";
        when "11111010110" => n11 <= "100000000100001111111101111100001001";
        when "11111010111" => n11 <= "100000000100000011111101111111010001";
        when "11111011000" => n11 <= "100000000011110110111110000010011010";
        when "11111011001" => n11 <= "100000000011101010111110000101100011";
        when "11111011010" => n11 <= "100000000011011110111110001000101011";
        when "11111011011" => n11 <= "100000000011010011111110001011110100";
        when "11111011100" => n11 <= "100000000011000111111110001110111101";
        when "11111011101" => n11 <= "100000000010111100111110010010000110";
        when "11111011110" => n11 <= "100000000010110010111110010101001110";
        when "11111011111" => n11 <= "100000000010100111111110011000010111";
        when "11111100000" => n11 <= "100000000010011101111110011011100000";
        when "11111100001" => n11 <= "100000000010010100111110011110101001";
        when "11111100010" => n11 <= "100000000010001010111110100001110010";
        when "11111100011" => n11 <= "100000000010000001111110100100111011";
        when "11111100100" => n11 <= "100000000001111000111110101000000011";
        when "11111100101" => n11 <= "100000000001110000111110101011001100";
        when "11111100110" => n11 <= "100000000001101000111110101110010101";
        when "11111100111" => n11 <= "100000000001100000111110110001011110";
        when "11111101000" => n11 <= "100000000001011000111110110100100111";
        when "11111101001" => n11 <= "100000000001010001111110110111110000";
        when "11111101010" => n11 <= "100000000001001010111110111010111001";
        when "11111101011" => n11 <= "100000000001000100111110111110000010";
        when "11111101100" => n11 <= "100000000000111101111111000001001011";
        when "11111101101" => n11 <= "100000000000110111111111000100010100";
        when "11111101110" => n11 <= "100000000000110001111111000111011101";
        when "11111101111" => n11 <= "100000000000101100111111001010100110";
        when "11111110000" => n11 <= "100000000000100111111111001101101111";
        when "11111110001" => n11 <= "100000000000100010111111010000111000";
        when "11111110010" => n11 <= "100000000000011110111111010100000001";
        when "11111110011" => n11 <= "100000000000011010111111010111001010";
        when "11111110100" => n11 <= "100000000000010110111111011010010011";
        when "11111110101" => n11 <= "100000000000010010111111011101011100";
        when "11111110110" => n11 <= "100000000000001111111111100000100101";
        when "11111110111" => n11 <= "100000000000001100111111100011101110";
        when "11111111000" => n11 <= "100000000000001001111111100110110111";
        when "11111111001" => n11 <= "100000000000000111111111101010000000";
        when "11111111010" => n11 <= "100000000000000101111111101101001001";
        when "11111111011" => n11 <= "100000000000000011111111110000010010";
        when "11111111100" => n11 <= "100000000000000010111111110011011011";
        when "11111111101" => n11 <= "100000000000000001111111110110100100";
        when "11111111110" => n11 <= "100000000000000000111111111001101101";
        when "11111111111" => n11 <= "100000000000000000111111111100110110";
        when others => n11 <= "XXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX";
      end case;
    end if;
  end if;
end process;
n12 <= n11(35 downto 35) &
  n11(34 downto 34) &
  n11(33 downto 33) &
  n11(32 downto 32) &
  n11(31 downto 31) &
  n11(30 downto 30) &
  n11(29 downto 29) &
  n11(28 downto 28) &
  n11(27 downto 27) &
  n11(26 downto 26) &
  n11(25 downto 25) &
  n11(24 downto 24) &
  n11(23 downto 23) &
  n11(22 downto 22) &
  n11(21 downto 21) &
  n11(20 downto 20) &
  n11(19 downto 19) &
  n11(18 downto 18);
n13 <= n11(17 downto 17) &
  n11(16 downto 16) &
  n11(15 downto 15) &
  n11(14 downto 14) &
  n11(13 downto 13) &
  n11(12 downto 12) &
  n11(11 downto 11) &
  n11(10 downto 10) &
  n11(9 downto 9) &
  n11(8 downto 8) &
  n11(7 downto 7) &
  n11(6 downto 6) &
  n11(5 downto 5) &
  n11(4 downto 4) &
  n11(3 downto 3) &
  n11(2 downto 2) &
  n11(1 downto 1) &
  n11(0 downto 0);
n14 <= unsigned(signed(n5) * signed(n12));
n15 <= n14(34 downto 34) &
  n14(33 downto 33) &
  n14(32 downto 32) &
  n14(31 downto 31) &
  n14(30 downto 30) &
  n14(29 downto 29) &
  n14(28 downto 28) &
  n14(27 downto 27) &
  n14(26 downto 26) &
  n14(25 downto 25) &
  n14(24 downto 24) &
  n14(23 downto 23) &
  n14(22 downto 22) &
  n14(21 downto 21) &
  n14(20 downto 20) &
  n14(19 downto 19) &
  n14(18 downto 18) &
  n14(17 downto 17);
process (clock_c) begin
  if rising_edge(clock_c) then
    if i5 = "1" then
      n16 <= "000000000000000000";
    elsif i4 = "1" then
      n16 <= n15;
    end if;
  end if;
end process;
n17 <= unsigned(signed(n6) * signed(n13));
n18 <= n17(34 downto 34) &
  n17(33 downto 33) &
  n17(32 downto 32) &
  n17(31 downto 31) &
  n17(30 downto 30) &
  n17(29 downto 29) &
  n17(28 downto 28) &
  n17(27 downto 27) &
  n17(26 downto 26) &
  n17(25 downto 25) &
  n17(24 downto 24) &
  n17(23 downto 23) &
  n17(22 downto 22) &
  n17(21 downto 21) &
  n17(20 downto 20) &
  n17(19 downto 19) &
  n17(18 downto 18) &
  n17(17 downto 17);
process (clock_c) begin
  if rising_edge(clock_c) then
    if i5 = "1" then
      n19 <= "000000000000000000";
    elsif i4 = "1" then
      n19 <= n18;
    end if;
  end if;
end process;
n20 <= n16 - n19;
process (clock_c) begin
  if rising_edge(clock_c) then
    if i5 = "1" then
      n21 <= "000000000000000000";
    elsif i4 = "1" then
      n21 <= n20;
    end if;
  end if;
end process;
n22 <= unsigned(signed(n5) * signed(n13));
n23 <= n22(34 downto 34) &
  n22(33 downto 33) &
  n22(32 downto 32) &
  n22(31 downto 31) &
  n22(30 downto 30) &
  n22(29 downto 29) &
  n22(28 downto 28) &
  n22(27 downto 27) &
  n22(26 downto 26) &
  n22(25 downto 25) &
  n22(24 downto 24) &
  n22(23 downto 23) &
  n22(22 downto 22) &
  n22(21 downto 21) &
  n22(20 downto 20) &
  n22(19 downto 19) &
  n22(18 downto 18) &
  n22(17 downto 17);
process (clock_c) begin
  if rising_edge(clock_c) then
    if i5 = "1" then
      n24 <= "000000000000000000";
    elsif i4 = "1" then
      n24 <= n23;
    end if;
  end if;
end process;
n25 <= unsigned(signed(n6) * signed(n12));
n26 <= n25(34 downto 34) &
  n25(33 downto 33) &
  n25(32 downto 32) &
  n25(31 downto 31) &
  n25(30 downto 30) &
  n25(29 downto 29) &
  n25(28 downto 28) &
  n25(27 downto 27) &
  n25(26 downto 26) &
  n25(25 downto 25) &
  n25(24 downto 24) &
  n25(23 downto 23) &
  n25(22 downto 22) &
  n25(21 downto 21) &
  n25(20 downto 20) &
  n25(19 downto 19) &
  n25(18 downto 18) &
  n25(17 downto 17);
process (clock_c) begin
  if rising_edge(clock_c) then
    if i5 = "1" then
      n27 <= "000000000000000000";
    elsif i4 = "1" then
      n27 <= n26;
    end if;
  end if;
end process;
n28 <= n24 + n27;
process (clock_c) begin
  if rising_edge(clock_c) then
    if i5 = "1" then
      n29 <= "000000000000000000";
    elsif i4 = "1" then
      n29 <= n28;
    end if;
  end if;
end process;
n30 <= n8 + n21;
n31 <= n10 + n29;
n32 <= n30 & n31;
process (clock_c) begin
  if rising_edge(clock_c) then
    if i5 = "1" then
      n33 <= "000000000000000000000000000000000000";
    elsif i4 = "1" then
      n33 <= n32;
    end if;
  end if;
end process;
n34 <= n8 - n21;
n35 <= n10 - n29;
n36 <= n34 & n35;
process (clock_c) begin
  if rising_edge(clock_c) then
    if i5 = "1" then
      n37 <= "000000000000000000000000000000000000";
    elsif i4 = "1" then
      n37 <= n36;
    end if;
  end if;
end process;
o2 <= n37;
o1 <= n33;
end architecture rtl;

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
entity cf_fft_4096_18_25 is
port (
clock_c : in std_logic;
i1 : in  unsigned(0 downto 0);
i2 : in  unsigned(35 downto 0);
i3 : in  unsigned(35 downto 0);
i4 : in  unsigned(0 downto 0);
i5 : in  unsigned(0 downto 0);
o1 : out unsigned(0 downto 0);
o2 : out unsigned(35 downto 0);
o3 : out unsigned(35 downto 0));
end entity cf_fft_4096_18_25;
architecture rtl of cf_fft_4096_18_25 is
signal n1 : unsigned(10 downto 0);
signal n2 : unsigned(71 downto 0);
signal n3 : unsigned(0 downto 0) := "0";
signal n4 : unsigned(0 downto 0) := "0";
signal n5 : unsigned(0 downto 0) := "0";
signal n6 : unsigned(0 downto 0) := "0";
signal n7 : unsigned(9 downto 0);
signal n8 : unsigned(9 downto 0) := "0000000000";
signal n9 : unsigned(9 downto 0) := "0000000000";
signal n10 : unsigned(9 downto 0) := "0000000000";
signal n11 : unsigned(9 downto 0) := "0000000000";
signal n12 : unsigned(0 downto 0);
signal n13 : unsigned(0 downto 0) := "0";
signal n14 : unsigned(0 downto 0) := "0";
signal n15 : unsigned(0 downto 0) := "0";
signal n16 : unsigned(0 downto 0) := "0";
signal n17 : unsigned(0 downto 0);
signal n18 : unsigned(1 downto 0);
signal n19 : unsigned(35 downto 0);
signal n20 : unsigned(35 downto 0);
signal n21 : unsigned(35 downto 0);
signal n22 : unsigned(35 downto 0);
signal n23 : unsigned(35 downto 0);
signal n24 : unsigned(35 downto 0);
signal s25_1 : unsigned(35 downto 0);
signal s25_2 : unsigned(35 downto 0);
signal s26_1 : unsigned(0 downto 0);
signal s27_1 : unsigned(71 downto 0);
signal s28_1 : unsigned(0 downto 0);
signal s28_2 : unsigned(0 downto 0);
signal s28_3 : unsigned(71 downto 0);
signal s29_1 : unsigned(10 downto 0);
signal s29_2 : unsigned(0 downto 0);
component cf_fft_4096_18_26 is
port (
clock_c : in std_logic;
i1 : in  unsigned(35 downto 0);
i2 : in  unsigned(35 downto 0);
i3 : in  unsigned(10 downto 0);
i4 : in  unsigned(0 downto 0);
i5 : in  unsigned(0 downto 0);
o1 : out unsigned(35 downto 0);
o2 : out unsigned(35 downto 0));
end component cf_fft_4096_18_26;
component cf_fft_4096_18_37 is
port (
clock_c : in std_logic;
i1 : in  unsigned(1 downto 0);
i2 : in  unsigned(0 downto 0);
i3 : in  unsigned(0 downto 0);
o1 : out unsigned(0 downto 0));
end component cf_fft_4096_18_37;
component cf_fft_4096_18_33 is
port (
clock_c : in std_logic;
i1 : in  unsigned(71 downto 0);
i2 : in  unsigned(0 downto 0);
i3 : in  unsigned(9 downto 0);
i4 : in  unsigned(0 downto 0);
i5 : in  unsigned(0 downto 0);
i6 : in  unsigned(0 downto 0);
o1 : out unsigned(71 downto 0));
end component cf_fft_4096_18_33;
component cf_fft_4096_18_32 is
port (
clock_c : in std_logic;
i1 : in  unsigned(71 downto 0);
i2 : in  unsigned(0 downto 0);
i3 : in  unsigned(9 downto 0);
i4 : in  unsigned(0 downto 0);
i5 : in  unsigned(0 downto 0);
i6 : in  unsigned(0 downto 0);
o1 : out unsigned(0 downto 0);
o2 : out unsigned(0 downto 0);
o3 : out unsigned(71 downto 0));
end component cf_fft_4096_18_32;
component cf_fft_4096_18_28 is
port (
clock_c : in std_logic;
i1 : in  unsigned(0 downto 0);
i2 : in  unsigned(0 downto 0);
i3 : in  unsigned(0 downto 0);
o1 : out unsigned(10 downto 0);
o2 : out unsigned(0 downto 0));
end component cf_fft_4096_18_28;
begin
n1 <= s29_1(10 downto 10) &
  s29_1(9 downto 9) &
  s29_1(8 downto 8) &
  s29_1(7 downto 7) &
  s29_1(6 downto 6) &
  s29_1(5 downto 5) &
  s29_1(4 downto 4) &
  s29_1(3 downto 3) &
  s29_1(2 downto 2) &
  s29_1(1 downto 1) &
  s29_1(0 downto 0);
n2 <= s25_1 & s25_2;
process (clock_c) begin
  if rising_edge(clock_c) then
    if i5 = "1" then
      n3 <= "0";
    elsif i4 = "1" then
      n3 <= s29_2;
    end if;
  end if;
end process;
process (clock_c) begin
  if rising_edge(clock_c) then
    if i5 = "1" then
      n4 <= "0";
    elsif i4 = "1" then
      n4 <= n3;
    end if;
  end if;
end process;
process (clock_c) begin
  if rising_edge(clock_c) then
    if i5 = "1" then
      n5 <= "0";
    elsif i4 = "1" then
      n5 <= n4;
    end if;
  end if;
end process;
process (clock_c) begin
  if rising_edge(clock_c) then
    if i5 = "1" then
      n6 <= "0";
    elsif i4 = "1" then
      n6 <= n5;
    end if;
  end if;
end process;
n7 <= s29_1(10 downto 10) &
  s29_1(9 downto 9) &
  s29_1(8 downto 8) &
  s29_1(7 downto 7) &
  s29_1(6 downto 6) &
  s29_1(5 downto 5) &
  s29_1(4 downto 4) &
  s29_1(3 downto 3) &
  s29_1(2 downto 2) &
  s29_1(1 downto 1);
process (clock_c) begin
  if rising_edge(clock_c) then
    if i5 = "1" then
      n8 <= "0000000000";
    elsif i4 = "1" then
      n8 <= n7;
    end if;
  end if;
end process;
process (clock_c) begin
  if rising_edge(clock_c) then
    if i5 = "1" then
      n9 <= "0000000000";
    elsif i4 = "1" then
      n9 <= n8;
    end if;
  end if;
end process;
process (clock_c) begin
  if rising_edge(clock_c) then
    if i5 = "1" then
      n10 <= "0000000000";
    elsif i4 = "1" then
      n10 <= n9;
    end if;
  end if;
end process;
process (clock_c) begin
  if rising_edge(clock_c) then
    if i5 = "1" then
      n11 <= "0000000000";
    elsif i4 = "1" then
      n11 <= n10;
    end if;
  end if;
end process;
n12 <= s29_1(0 downto 0);
process (clock_c) begin
  if rising_edge(clock_c) then
    if i5 = "1" then
      n13 <= "0";
    elsif i4 = "1" then
      n13 <= n12;
    end if;
  end if;
end process;
process (clock_c) begin
  if rising_edge(clock_c) then
    if i5 = "1" then
      n14 <= "0";
    elsif i4 = "1" then
      n14 <= n13;
    end if;
  end if;
end process;
process (clock_c) begin
  if rising_edge(clock_c) then
    if i5 = "1" then
      n15 <= "0";
    elsif i4 = "1" then
      n15 <= n14;
    end if;
  end if;
end process;
process (clock_c) begin
  if rising_edge(clock_c) then
    if i5 = "1" then
      n16 <= "0";
    elsif i4 = "1" then
      n16 <= n15;
    end if;
  end if;
end process;
n17 <= not n16;
n18 <= s28_2 & s28_1;
n19 <= s28_3(71 downto 71) &
  s28_3(70 downto 70) &
  s28_3(69 downto 69) &
  s28_3(68 downto 68) &
  s28_3(67 downto 67) &
  s28_3(66 downto 66) &
  s28_3(65 downto 65) &
  s28_3(64 downto 64) &
  s28_3(63 downto 63) &
  s28_3(62 downto 62) &
  s28_3(61 downto 61) &
  s28_3(60 downto 60) &
  s28_3(59 downto 59) &
  s28_3(58 downto 58) &
  s28_3(57 downto 57) &
  s28_3(56 downto 56) &
  s28_3(55 downto 55) &
  s28_3(54 downto 54) &
  s28_3(53 downto 53) &
  s28_3(52 downto 52) &
  s28_3(51 downto 51) &
  s28_3(50 downto 50) &
  s28_3(49 downto 49) &
  s28_3(48 downto 48) &
  s28_3(47 downto 47) &
  s28_3(46 downto 46) &
  s28_3(45 downto 45) &
  s28_3(44 downto 44) &
  s28_3(43 downto 43) &
  s28_3(42 downto 42) &
  s28_3(41 downto 41) &
  s28_3(40 downto 40) &
  s28_3(39 downto 39) &
  s28_3(38 downto 38) &
  s28_3(37 downto 37) &
  s28_3(36 downto 36);
n20 <= s28_3(35 downto 35) &
  s28_3(34 downto 34) &
  s28_3(33 downto 33) &
  s28_3(32 downto 32) &
  s28_3(31 downto 31) &
  s28_3(30 downto 30) &
  s28_3(29 downto 29) &
  s28_3(28 downto 28) &
  s28_3(27 downto 27) &
  s28_3(26 downto 26) &
  s28_3(25 downto 25) &
  s28_3(24 downto 24) &
  s28_3(23 downto 23) &
  s28_3(22 downto 22) &
  s28_3(21 downto 21) &
  s28_3(20 downto 20) &
  s28_3(19 downto 19) &
  s28_3(18 downto 18) &
  s28_3(17 downto 17) &
  s28_3(16 downto 16) &
  s28_3(15 downto 15) &
  s28_3(14 downto 14) &
  s28_3(13 downto 13) &
  s28_3(12 downto 12) &
  s28_3(11 downto 11) &
  s28_3(10 downto 10) &
  s28_3(9 downto 9) &
  s28_3(8 downto 8) &
  s28_3(7 downto 7) &
  s28_3(6 downto 6) &
  s28_3(5 downto 5) &
  s28_3(4 downto 4) &
  s28_3(3 downto 3) &
  s28_3(2 downto 2) &
  s28_3(1 downto 1) &
  s28_3(0 downto 0);
n21 <= s27_1(71 downto 71) &
  s27_1(70 downto 70) &
  s27_1(69 downto 69) &
  s27_1(68 downto 68) &
  s27_1(67 downto 67) &
  s27_1(66 downto 66) &
  s27_1(65 downto 65) &
  s27_1(64 downto 64) &
  s27_1(63 downto 63) &
  s27_1(62 downto 62) &
  s27_1(61 downto 61) &
  s27_1(60 downto 60) &
  s27_1(59 downto 59) &
  s27_1(58 downto 58) &
  s27_1(57 downto 57) &
  s27_1(56 downto 56) &
  s27_1(55 downto 55) &
  s27_1(54 downto 54) &
  s27_1(53 downto 53) &
  s27_1(52 downto 52) &
  s27_1(51 downto 51) &
  s27_1(50 downto 50) &
  s27_1(49 downto 49) &
  s27_1(48 downto 48) &
  s27_1(47 downto 47) &
  s27_1(46 downto 46) &
  s27_1(45 downto 45) &
  s27_1(44 downto 44) &
  s27_1(43 downto 43) &
  s27_1(42 downto 42) &
  s27_1(41 downto 41) &
  s27_1(40 downto 40) &
  s27_1(39 downto 39) &
  s27_1(38 downto 38) &
  s27_1(37 downto 37) &
  s27_1(36 downto 36);
n22 <= s27_1(35 downto 35) &
  s27_1(34 downto 34) &
  s27_1(33 downto 33) &
  s27_1(32 downto 32) &
  s27_1(31 downto 31) &
  s27_1(30 downto 30) &
  s27_1(29 downto 29) &
  s27_1(28 downto 28) &
  s27_1(27 downto 27) &
  s27_1(26 downto 26) &
  s27_1(25 downto 25) &
  s27_1(24 downto 24) &
  s27_1(23 downto 23) &
  s27_1(22 downto 22) &
  s27_1(21 downto 21) &
  s27_1(20 downto 20) &
  s27_1(19 downto 19) &
  s27_1(18 downto 18) &
  s27_1(17 downto 17) &
  s27_1(16 downto 16) &
  s27_1(15 downto 15) &
  s27_1(14 downto 14) &
  s27_1(13 downto 13) &
  s27_1(12 downto 12) &
  s27_1(11 downto 11) &
  s27_1(10 downto 10) &
  s27_1(9 downto 9) &
  s27_1(8 downto 8) &
  s27_1(7 downto 7) &
  s27_1(6 downto 6) &
  s27_1(5 downto 5) &
  s27_1(4 downto 4) &
  s27_1(3 downto 3) &
  s27_1(2 downto 2) &
  s27_1(1 downto 1) &
  s27_1(0 downto 0);
n23 <= n20 when s26_1 = "1" else n19;
n24 <= n22 when s26_1 = "1" else n21;
s25 : cf_fft_4096_18_26 port map (clock_c, i2, i3, n1, i4, i5, s25_1, s25_2);
s26 : cf_fft_4096_18_37 port map (clock_c, n18, i4, i5, s26_1);
s27 : cf_fft_4096_18_33 port map (clock_c, n2, n6, n11, n16, i4, i5, s27_1);
s28 : cf_fft_4096_18_32 port map (clock_c, n2, n6, n11, n17, i4, i5, s28_1, s28_2, s28_3);
s29 : cf_fft_4096_18_28 port map (clock_c, i1, i4, i5, s29_1, s29_2);
o3 <= n24;
o2 <= n23;
o1 <= s28_1;
end architecture rtl;

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
entity cf_fft_4096_18_24 is
port (
clock_c : in std_logic;
i1 : in  unsigned(35 downto 0);
i2 : in  unsigned(35 downto 0);
i3 : in  unsigned(9 downto 0);
i4 : in  unsigned(0 downto 0);
i5 : in  unsigned(0 downto 0);
o1 : out unsigned(35 downto 0);
o2 : out unsigned(35 downto 0));
end entity cf_fft_4096_18_24;
architecture rtl of cf_fft_4096_18_24 is
signal n1 : unsigned(35 downto 0) := "000000000000000000000000000000000000";
signal n2 : unsigned(17 downto 0);
signal n3 : unsigned(17 downto 0);
signal n4 : unsigned(35 downto 0) := "000000000000000000000000000000000000";
signal n5 : unsigned(17 downto 0);
signal n6 : unsigned(17 downto 0);
signal n7 : unsigned(17 downto 0) := "000000000000000000";
signal n8 : unsigned(17 downto 0) := "000000000000000000";
signal n9 : unsigned(17 downto 0) := "000000000000000000";
signal n10 : unsigned(17 downto 0) := "000000000000000000";
signal n11 : unsigned(35 downto 0) := "000000000000000000000000000000000000";
signal n12 : unsigned(17 downto 0);
signal n13 : unsigned(17 downto 0);
signal n14 : unsigned(35 downto 0);
signal n15 : unsigned(17 downto 0);
signal n16 : unsigned(17 downto 0) := "000000000000000000";
signal n17 : unsigned(35 downto 0);
signal n18 : unsigned(17 downto 0);
signal n19 : unsigned(17 downto 0) := "000000000000000000";
signal n20 : unsigned(17 downto 0);
signal n21 : unsigned(17 downto 0) := "000000000000000000";
signal n22 : unsigned(35 downto 0);
signal n23 : unsigned(17 downto 0);
signal n24 : unsigned(17 downto 0) := "000000000000000000";
signal n25 : unsigned(35 downto 0);
signal n26 : unsigned(17 downto 0);
signal n27 : unsigned(17 downto 0) := "000000000000000000";
signal n28 : unsigned(17 downto 0);
signal n29 : unsigned(17 downto 0) := "000000000000000000";
signal n30 : unsigned(17 downto 0);
signal n31 : unsigned(17 downto 0);
signal n32 : unsigned(35 downto 0);
signal n33 : unsigned(35 downto 0) := "000000000000000000000000000000000000";
signal n34 : unsigned(17 downto 0);
signal n35 : unsigned(17 downto 0);
signal n36 : unsigned(35 downto 0);
signal n37 : unsigned(35 downto 0) := "000000000000000000000000000000000000";
begin
process (clock_c) begin
  if rising_edge(clock_c) then
    if i5 = "1" then
      n1 <= "000000000000000000000000000000000000";
    elsif i4 = "1" then
      n1 <= i1;
    end if;
  end if;
end process;
n2 <= n1(35 downto 35) &
  n1(34 downto 34) &
  n1(33 downto 33) &
  n1(32 downto 32) &
  n1(31 downto 31) &
  n1(30 downto 30) &
  n1(29 downto 29) &
  n1(28 downto 28) &
  n1(27 downto 27) &
  n1(26 downto 26) &
  n1(25 downto 25) &
  n1(24 downto 24) &
  n1(23 downto 23) &
  n1(22 downto 22) &
  n1(21 downto 21) &
  n1(20 downto 20) &
  n1(19 downto 19) &
  n1(18 downto 18);
n3 <= n1(17 downto 17) &
  n1(16 downto 16) &
  n1(15 downto 15) &
  n1(14 downto 14) &
  n1(13 downto 13) &
  n1(12 downto 12) &
  n1(11 downto 11) &
  n1(10 downto 10) &
  n1(9 downto 9) &
  n1(8 downto 8) &
  n1(7 downto 7) &
  n1(6 downto 6) &
  n1(5 downto 5) &
  n1(4 downto 4) &
  n1(3 downto 3) &
  n1(2 downto 2) &
  n1(1 downto 1) &
  n1(0 downto 0);
process (clock_c) begin
  if rising_edge(clock_c) then
    if i5 = "1" then
      n4 <= "000000000000000000000000000000000000";
    elsif i4 = "1" then
      n4 <= i2;
    end if;
  end if;
end process;
n5 <= n4(35 downto 35) &
  n4(34 downto 34) &
  n4(33 downto 33) &
  n4(32 downto 32) &
  n4(31 downto 31) &
  n4(30 downto 30) &
  n4(29 downto 29) &
  n4(28 downto 28) &
  n4(27 downto 27) &
  n4(26 downto 26) &
  n4(25 downto 25) &
  n4(24 downto 24) &
  n4(23 downto 23) &
  n4(22 downto 22) &
  n4(21 downto 21) &
  n4(20 downto 20) &
  n4(19 downto 19) &
  n4(18 downto 18);
n6 <= n4(17 downto 17) &
  n4(16 downto 16) &
  n4(15 downto 15) &
  n4(14 downto 14) &
  n4(13 downto 13) &
  n4(12 downto 12) &
  n4(11 downto 11) &
  n4(10 downto 10) &
  n4(9 downto 9) &
  n4(8 downto 8) &
  n4(7 downto 7) &
  n4(6 downto 6) &
  n4(5 downto 5) &
  n4(4 downto 4) &
  n4(3 downto 3) &
  n4(2 downto 2) &
  n4(1 downto 1) &
  n4(0 downto 0);
process (clock_c) begin
  if rising_edge(clock_c) then
    if i5 = "1" then
      n7 <= "000000000000000000";
    elsif i4 = "1" then
      n7 <= n2;
    end if;
  end if;
end process;
process (clock_c) begin
  if rising_edge(clock_c) then
    if i5 = "1" then
      n8 <= "000000000000000000";
    elsif i4 = "1" then
      n8 <= n7;
    end if;
  end if;
end process;
process (clock_c) begin
  if rising_edge(clock_c) then
    if i5 = "1" then
      n9 <= "000000000000000000";
    elsif i4 = "1" then
      n9 <= n3;
    end if;
  end if;
end process;
process (clock_c) begin
  if rising_edge(clock_c) then
    if i5 = "1" then
      n10 <= "000000000000000000";
    elsif i4 = "1" then
      n10 <= n9;
    end if;
  end if;
end process;
process (clock_c) begin
  if rising_edge(clock_c) then 
    if i4 = "1" then
      case i3 is
        when "0000000000" => n11 <= "011111111111111111000000000000000000";
        when "0000000001" => n11 <= "011111111111111111111111111001101101";
        when "0000000010" => n11 <= "011111111111111101111111110011011011";
        when "0000000011" => n11 <= "011111111111111010111111101101001001";
        when "0000000100" => n11 <= "011111111111110110111111100110110111";
        when "0000000101" => n11 <= "011111111111110000111111100000100101";
        when "0000000110" => n11 <= "011111111111101001111111011010010011";
        when "0000000111" => n11 <= "011111111111100001111111010100000001";
        when "0000001000" => n11 <= "011111111111011000111111001101101111";
        when "0000001001" => n11 <= "011111111111001110111111000111011101";
        when "0000001010" => n11 <= "011111111111000010111111000001001011";
        when "0000001011" => n11 <= "011111111110110101111110111010111001";
        when "0000001100" => n11 <= "011111111110100111111110110100100111";
        when "0000001101" => n11 <= "011111111110010111111110101110010101";
        when "0000001110" => n11 <= "011111111110000111111110101000000011";
        when "0000001111" => n11 <= "011111111101110101111110100001110010";
        when "0000010000" => n11 <= "011111111101100010111110011011100000";
        when "0000010001" => n11 <= "011111111101001101111110010101001110";
        when "0000010010" => n11 <= "011111111100111000111110001110111101";
        when "0000010011" => n11 <= "011111111100100001111110001000101011";
        when "0000010100" => n11 <= "011111111100001001111110000010011010";
        when "0000010101" => n11 <= "011111111011110000111101111100001001";
        when "0000010110" => n11 <= "011111111011010101111101110101110111";
        when "0000010111" => n11 <= "011111111010111001111101101111100110";
        when "0000011000" => n11 <= "011111111010011100111101101001010101";
        when "0000011001" => n11 <= "011111111001111110111101100011000100";
        when "0000011010" => n11 <= "011111111001011111111101011100110011";
        when "0000011011" => n11 <= "011111111000111110111101010110100011";
        when "0000011100" => n11 <= "011111111000011100111101010000010010";
        when "0000011101" => n11 <= "011111110111111001111101001010000001";
        when "0000011110" => n11 <= "011111110111010101111101000011110001";
        when "0000011111" => n11 <= "011111110110101111111100111101100000";
        when "0000100000" => n11 <= "011111110110001000111100110111010000";
        when "0000100001" => n11 <= "011111110101100000111100110001000000";
        when "0000100010" => n11 <= "011111110100110111111100101010110000";
        when "0000100011" => n11 <= "011111110100001101111100100100100000";
        when "0000100100" => n11 <= "011111110011100001111100011110010000";
        when "0000100101" => n11 <= "011111110010110100111100011000000001";
        when "0000100110" => n11 <= "011111110010000110111100010001110001";
        when "0000100111" => n11 <= "011111110001010110111100001011100010";
        when "0000101000" => n11 <= "011111110000100110111100000101010011";
        when "0000101001" => n11 <= "011111101111110100111011111111000100";
        when "0000101010" => n11 <= "011111101111000001111011111000110101";
        when "0000101011" => n11 <= "011111101110001101111011110010100110";
        when "0000101100" => n11 <= "011111101101010111111011101100011000";
        when "0000101101" => n11 <= "011111101100100000111011100110001001";
        when "0000101110" => n11 <= "011111101011101000111011011111111011";
        when "0000101111" => n11 <= "011111101010101111111011011001101101";
        when "0000110000" => n11 <= "011111101001110101111011010011011111";
        when "0000110001" => n11 <= "011111101000111001111011001101010010";
        when "0000110010" => n11 <= "011111100111111100111011000111000100";
        when "0000110011" => n11 <= "011111100110111110111011000000110111";
        when "0000110100" => n11 <= "011111100101111111111010111010101010";
        when "0000110101" => n11 <= "011111100100111111111010110100011101";
        when "0000110110" => n11 <= "011111100011111101111010101110010000";
        when "0000110111" => n11 <= "011111100010111010111010101000000011";
        when "0000111000" => n11 <= "011111100001110110111010100001110111";
        when "0000111001" => n11 <= "011111100000110000111010011011101011";
        when "0000111010" => n11 <= "011111011111101010111010010101011111";
        when "0000111011" => n11 <= "011111011110100010111010001111010100";
        when "0000111100" => n11 <= "011111011101011001111010001001001000";
        when "0000111101" => n11 <= "011111011100001111111010000010111101";
        when "0000111110" => n11 <= "011111011011000011111001111100110010";
        when "0000111111" => n11 <= "011111011001110111111001110110100111";
        when "0001000000" => n11 <= "011111011000101001111001110000011101";
        when "0001000001" => n11 <= "011111010111011010111001101010010010";
        when "0001000010" => n11 <= "011111010110001010111001100100001000";
        when "0001000011" => n11 <= "011111010100111000111001011101111111";
        when "0001000100" => n11 <= "011111010011100110111001010111110101";
        when "0001000101" => n11 <= "011111010010010010111001010001101100";
        when "0001000110" => n11 <= "011111010000111101111001001011100011";
        when "0001000111" => n11 <= "011111001111100110111001000101011010";
        when "0001001000" => n11 <= "011111001110001111111000111111010001";
        when "0001001001" => n11 <= "011111001100110110111000111001001001";
        when "0001001010" => n11 <= "011111001011011100111000110011000001";
        when "0001001011" => n11 <= "011111001010000001111000101100111010";
        when "0001001100" => n11 <= "011111001000100101111000100110110010";
        when "0001001101" => n11 <= "011111000111000111111000100000101011";
        when "0001001110" => n11 <= "011111000101101000111000011010100100";
        when "0001001111" => n11 <= "011111000100001001111000010100011110";
        when "0001010000" => n11 <= "011111000010100111111000001110011000";
        when "0001010001" => n11 <= "011111000001000101111000001000010010";
        when "0001010010" => n11 <= "011110111111100010111000000010001100";
        when "0001010011" => n11 <= "011110111101111101110111111100000111";
        when "0001010100" => n11 <= "011110111100010111110111110110000010";
        when "0001010101" => n11 <= "011110111010110000110111101111111101";
        when "0001010110" => n11 <= "011110111001001000110111101001111001";
        when "0001010111" => n11 <= "011110110111011110110111100011110101";
        when "0001011000" => n11 <= "011110110101110100110111011101110001";
        when "0001011001" => n11 <= "011110110100001000110111010111101110";
        when "0001011010" => n11 <= "011110110010011011110111010001101010";
        when "0001011011" => n11 <= "011110110000101100110111001011101000";
        when "0001011100" => n11 <= "011110101110111101110111000101100101";
        when "0001011101" => n11 <= "011110101101001100110110111111100011";
        when "0001011110" => n11 <= "011110101011011011110110111001100010";
        when "0001011111" => n11 <= "011110101001101000110110110011100000";
        when "0001100000" => n11 <= "011110100111110100110110101101011111";
        when "0001100001" => n11 <= "011110100101111110110110100111011111";
        when "0001100010" => n11 <= "011110100100001000110110100001011110";
        when "0001100011" => n11 <= "011110100010010000110110011011011111";
        when "0001100100" => n11 <= "011110100000010111110110010101011111";
        when "0001100101" => n11 <= "011110011110011101110110001111100000";
        when "0001100110" => n11 <= "011110011100100010110110001001100001";
        when "0001100111" => n11 <= "011110011010100110110110000011100011";
        when "0001101000" => n11 <= "011110011000101000110101111101100101";
        when "0001101001" => n11 <= "011110010110101001110101110111100111";
        when "0001101010" => n11 <= "011110010100101001110101110001101010";
        when "0001101011" => n11 <= "011110010010101000110101101011101101";
        when "0001101100" => n11 <= "011110010000100110110101100101110000";
        when "0001101101" => n11 <= "011110001110100011110101011111110100";
        when "0001101110" => n11 <= "011110001100011110110101011001111001";
        when "0001101111" => n11 <= "011110001010011000110101010011111101";
        when "0001110000" => n11 <= "011110001000010010110101001110000011";
        when "0001110001" => n11 <= "011110000110001010110101001000001000";
        when "0001110010" => n11 <= "011110000100000000110101000010001110";
        when "0001110011" => n11 <= "011110000001110110110100111100010101";
        when "0001110100" => n11 <= "011101111111101010110100110110011100";
        when "0001110101" => n11 <= "011101111101011110110100110000100011";
        when "0001110110" => n11 <= "011101111011010000110100101010101011";
        when "0001110111" => n11 <= "011101111001000001110100100100110011";
        when "0001111000" => n11 <= "011101110110110001110100011110111011";
        when "0001111001" => n11 <= "011101110100011111110100011001000100";
        when "0001111010" => n11 <= "011101110010001101110100010011001110";
        when "0001111011" => n11 <= "011101101111111001110100001101011000";
        when "0001111100" => n11 <= "011101101101100101110100000111100010";
        when "0001111101" => n11 <= "011101101011001111110100000001101101";
        when "0001111110" => n11 <= "011101101000111000110011111011111000";
        when "0001111111" => n11 <= "011101100110100000110011110110000100";
        when "0010000000" => n11 <= "011101100100000110110011110000010000";
        when "0010000001" => n11 <= "011101100001101100110011101010011101";
        when "0010000010" => n11 <= "011101011111010000110011100100101010";
        when "0010000011" => n11 <= "011101011100110011110011011110111000";
        when "0010000100" => n11 <= "011101011010010110110011011001000110";
        when "0010000101" => n11 <= "011101010111110111110011010011010101";
        when "0010000110" => n11 <= "011101010101010110110011001101100100";
        when "0010000111" => n11 <= "011101010010110101110011000111110100";
        when "0010001000" => n11 <= "011101010000010011110011000010000100";
        when "0010001001" => n11 <= "011101001101101111110010111100010100";
        when "0010001010" => n11 <= "011101001011001011110010110110100101";
        when "0010001011" => n11 <= "011101001000100101110010110000110111";
        when "0010001100" => n11 <= "011101000101111110110010101011001001";
        when "0010001101" => n11 <= "011101000011010110110010100101011100";
        when "0010001110" => n11 <= "011101000000101101110010011111101111";
        when "0010001111" => n11 <= "011100111110000011110010011010000011";
        when "0010010000" => n11 <= "011100111011010111110010010100010111";
        when "0010010001" => n11 <= "011100111000101011110010001110101100";
        when "0010010010" => n11 <= "011100110101111101110010001001000001";
        when "0010010011" => n11 <= "011100110011001110110010000011010111";
        when "0010010100" => n11 <= "011100110000011111110001111101101101";
        when "0010010101" => n11 <= "011100101101101110110001111000000100";
        when "0010010110" => n11 <= "011100101010111100110001110010011100";
        when "0010010111" => n11 <= "011100101000001000110001101100110100";
        when "0010011000" => n11 <= "011100100101010100110001100111001100";
        when "0010011001" => n11 <= "011100100010011111110001100001100101";
        when "0010011010" => n11 <= "011100011111101000110001011011111111";
        when "0010011011" => n11 <= "011100011100110001110001010110011001";
        when "0010011100" => n11 <= "011100011001111000110001010000110100";
        when "0010011101" => n11 <= "011100010110111110110001001011001111";
        when "0010011110" => n11 <= "011100010100000100110001000101101011";
        when "0010011111" => n11 <= "011100010001001000110001000000001000";
        when "0010100000" => n11 <= "011100001110001011110000111010100101";
        when "0010100001" => n11 <= "011100001011001101110000110101000010";
        when "0010100010" => n11 <= "011100001000001101110000101111100000";
        when "0010100011" => n11 <= "011100000101001101110000101001111111";
        when "0010100100" => n11 <= "011100000010001100110000100100011111";
        when "0010100101" => n11 <= "011011111111001001110000011110111111";
        when "0010100110" => n11 <= "011011111100000110110000011001011111";
        when "0010100111" => n11 <= "011011111001000001110000010100000001";
        when "0010101000" => n11 <= "011011110101111100110000001110100010";
        when "0010101001" => n11 <= "011011110010110101110000001001000101";
        when "0010101010" => n11 <= "011011101111101101110000000011101000";
        when "0010101011" => n11 <= "011011101100100100101111111110001011";
        when "0010101100" => n11 <= "011011101001011010101111111000110000";
        when "0010101101" => n11 <= "011011100110001111101111110011010101";
        when "0010101110" => n11 <= "011011100011000011101111101101111010";
        when "0010101111" => n11 <= "011011011111110110101111101000100000";
        when "0010110000" => n11 <= "011011011100101000101111100011000111";
        when "0010110001" => n11 <= "011011011001011000101111011101101110";
        when "0010110010" => n11 <= "011011010110001000101111011000010110";
        when "0010110011" => n11 <= "011011010010110111101111010010111111";
        when "0010110100" => n11 <= "011011001111100100101111001101101000";
        when "0010110101" => n11 <= "011011001100010001101111001000010010";
        when "0010110110" => n11 <= "011011001000111100101111000010111101";
        when "0010110111" => n11 <= "011011000101100111101110111101101000";
        when "0010111000" => n11 <= "011011000010010000101110111000010100";
        when "0010111001" => n11 <= "011010111110111000101110110011000001";
        when "0010111010" => n11 <= "011010111011100000101110101101101110";
        when "0010111011" => n11 <= "011010111000000110101110101000011100";
        when "0010111100" => n11 <= "011010110100101011101110100011001011";
        when "0010111101" => n11 <= "011010110001001111101110011101111010";
        when "0010111110" => n11 <= "011010101101110011101110011000101010";
        when "0010111111" => n11 <= "011010101010010101101110010011011010";
        when "0011000000" => n11 <= "011010100110110110101110001110001100";
        when "0011000001" => n11 <= "011010100011010110101110001000111110";
        when "0011000010" => n11 <= "011010011111110101101110000011110000";
        when "0011000011" => n11 <= "011010011100010011101101111110100100";
        when "0011000100" => n11 <= "011010011000110000101101111001011000";
        when "0011000101" => n11 <= "011010010101001100101101110100001101";
        when "0011000110" => n11 <= "011010010001100111101101101111000010";
        when "0011000111" => n11 <= "011010001110000001101101101001111000";
        when "0011001000" => n11 <= "011010001010011010101101100100101111";
        when "0011001001" => n11 <= "011010000110110010101101011111100111";
        when "0011001010" => n11 <= "011010000011001001101101011010011111";
        when "0011001011" => n11 <= "011001111111011111101101010101011000";
        when "0011001100" => n11 <= "011001111011110100101101010000010010";
        when "0011001101" => n11 <= "011001111000001000101101001011001100";
        when "0011001110" => n11 <= "011001110100011011101101000110000111";
        when "0011001111" => n11 <= "011001110000101101101101000001000011";
        when "0011010000" => n11 <= "011001101100111110101100111100000000";
        when "0011010001" => n11 <= "011001101001001101101100110110111101";
        when "0011010010" => n11 <= "011001100101011100101100110001111011";
        when "0011010011" => n11 <= "011001100001101010101100101100111010";
        when "0011010100" => n11 <= "011001011101110111101100100111111010";
        when "0011010101" => n11 <= "011001011010000011101100100010111010";
        when "0011010110" => n11 <= "011001010110001110101100011101111011";
        when "0011010111" => n11 <= "011001010010011001101100011000111101";
        when "0011011000" => n11 <= "011001001110100010101100010100000000";
        when "0011011001" => n11 <= "011001001010101010101100001111000011";
        when "0011011010" => n11 <= "011001000110110001101100001010000111";
        when "0011011011" => n11 <= "011001000010110111101100000101001100";
        when "0011011100" => n11 <= "011000111110111100101100000000010010";
        when "0011011101" => n11 <= "011000111011000001101011111011011000";
        when "0011011110" => n11 <= "011000110111000100101011110110100000";
        when "0011011111" => n11 <= "011000110011000110101011110001101000";
        when "0011100000" => n11 <= "011000101111001000101011101100110000";
        when "0011100001" => n11 <= "011000101011001000101011100111111010";
        when "0011100010" => n11 <= "011000100111000111101011100011000100";
        when "0011100011" => n11 <= "011000100011000110101011011110001111";
        when "0011100100" => n11 <= "011000011111000100101011011001011011";
        when "0011100101" => n11 <= "011000011011000000101011010100101000";
        when "0011100110" => n11 <= "011000010110111100101011001111110101";
        when "0011100111" => n11 <= "011000010010110111101011001011000100";
        when "0011101000" => n11 <= "011000001110110000101011000110010011";
        when "0011101001" => n11 <= "011000001010101001101011000001100011";
        when "0011101010" => n11 <= "011000000110100001101010111100110011";
        when "0011101011" => n11 <= "011000000010011000101010111000000101";
        when "0011101100" => n11 <= "010111111110001110101010110011010111";
        when "0011101101" => n11 <= "010111111010000011101010101110101011";
        when "0011101110" => n11 <= "010111110101111000101010101001111110";
        when "0011101111" => n11 <= "010111110001101011101010100101010011";
        when "0011110000" => n11 <= "010111101101011101101010100000101001";
        when "0011110001" => n11 <= "010111101001001111101010011011111111";
        when "0011110010" => n11 <= "010111100101000000101010010111010111";
        when "0011110011" => n11 <= "010111100000101111101010010010101111";
        when "0011110100" => n11 <= "010111011100011110101010001110001000";
        when "0011110101" => n11 <= "010111011000001100101010001001100010";
        when "0011110110" => n11 <= "010111010011111001101010000100111100";
        when "0011110111" => n11 <= "010111001111100101101010000000011000";
        when "0011111000" => n11 <= "010111001011010000101001111011110100";
        when "0011111001" => n11 <= "010111000110111010101001110111010001";
        when "0011111010" => n11 <= "010111000010100100101001110010101111";
        when "0011111011" => n11 <= "010110111110001100101001101110001110";
        when "0011111100" => n11 <= "010110111001110100101001101001101110";
        when "0011111101" => n11 <= "010110110101011010101001100101001111";
        when "0011111110" => n11 <= "010110110001000000101001100000110000";
        when "0011111111" => n11 <= "010110101100100101101001011100010010";
        when "0100000000" => n11 <= "010110101000001001101001010111110110";
        when "0100000001" => n11 <= "010110100011101101101001010011011010";
        when "0100000010" => n11 <= "010110011111001111101001001110111111";
        when "0100000011" => n11 <= "010110011010110000101001001010100101";
        when "0100000100" => n11 <= "010110010110010001101001000110001011";
        when "0100000101" => n11 <= "010110010001110001101001000001110011";
        when "0100000110" => n11 <= "010110001101010000101000111101011011";
        when "0100000111" => n11 <= "010110001000101110101000111001000101";
        when "0100001000" => n11 <= "010110000100001011101000110100101111";
        when "0100001001" => n11 <= "010101111111100111101000110000011010";
        when "0100001010" => n11 <= "010101111011000011101000101100000110";
        when "0100001011" => n11 <= "010101110110011101101000100111110011";
        when "0100001100" => n11 <= "010101110001110111101000100011100001";
        when "0100001101" => n11 <= "010101101101010000101000011111010000";
        when "0100001110" => n11 <= "010101101000101000101000011010111111";
        when "0100001111" => n11 <= "010101100100000000101000010110110000";
        when "0100010000" => n11 <= "010101011111010110101000010010100010";
        when "0100010001" => n11 <= "010101011010101100101000001110010100";
        when "0100010010" => n11 <= "010101010110000001101000001010000111";
        when "0100010011" => n11 <= "010101010001010100101000000101111100";
        when "0100010100" => n11 <= "010101001100101000101000000001110001";
        when "0100010101" => n11 <= "010101000111111010100111111101100111";
        when "0100010110" => n11 <= "010101000011001100100111111001011110";
        when "0100010111" => n11 <= "010100111110011100100111110101010110";
        when "0100011000" => n11 <= "010100111001101100100111110001001111";
        when "0100011001" => n11 <= "010100110100111011100111101101001000";
        when "0100011010" => n11 <= "010100110000001010100111101001000011";
        when "0100011011" => n11 <= "010100101011010111100111100100111111";
        when "0100011100" => n11 <= "010100100110100100100111100000111011";
        when "0100011101" => n11 <= "010100100001110000100111011100111001";
        when "0100011110" => n11 <= "010100011100111011100111011000111000";
        when "0100011111" => n11 <= "010100011000000101100111010100110111";
        when "0100100000" => n11 <= "010100010011001111100111010000110111";
        when "0100100001" => n11 <= "010100001110010111100111001100111001";
        when "0100100010" => n11 <= "010100001001011111100111001000111011";
        when "0100100011" => n11 <= "010100000100100111100111000100111110";
        when "0100100100" => n11 <= "010011111111101101100111000001000011";
        when "0100100101" => n11 <= "010011111010110011100110111101001000";
        when "0100100110" => n11 <= "010011110101111000100110111001001110";
        when "0100100111" => n11 <= "010011110000111100100110110101010101";
        when "0100101000" => n11 <= "010011101011111111100110110001011101";
        when "0100101001" => n11 <= "010011100111000010100110101101100110";
        when "0100101010" => n11 <= "010011100010000100100110101001110001";
        when "0100101011" => n11 <= "010011011101000101100110100101111100";
        when "0100101100" => n11 <= "010011011000000101100110100010001000";
        when "0100101101" => n11 <= "010011010011000101100110011110010101";
        when "0100101110" => n11 <= "010011001110000100100110011010100011";
        when "0100101111" => n11 <= "010011001001000010100110010110110010";
        when "0100110000" => n11 <= "010011000011111111100110010011000001";
        when "0100110001" => n11 <= "010010111110111100100110001111010010";
        when "0100110010" => n11 <= "010010111001111000100110001011100100";
        when "0100110011" => n11 <= "010010110100110011100110000111110111";
        when "0100110100" => n11 <= "010010101111101101100110000100001011";
        when "0100110101" => n11 <= "010010101010100111100110000000100000";
        when "0100110110" => n11 <= "010010100101100000100101111100110110";
        when "0100110111" => n11 <= "010010100000011000100101111001001101";
        when "0100111000" => n11 <= "010010011011010000100101110101100101";
        when "0100111001" => n11 <= "010010010110000111100101110001111110";
        when "0100111010" => n11 <= "010010010000111101100101101110011000";
        when "0100111011" => n11 <= "010010001011110010100101101010110011";
        when "0100111100" => n11 <= "010010000110100111100101100111001111";
        when "0100111101" => n11 <= "010010000001011011100101100011101100";
        when "0100111110" => n11 <= "010001111100001111100101100000001010";
        when "0100111111" => n11 <= "010001110111000001100101011100101001";
        when "0101000000" => n11 <= "010001110001110011100101011001001001";
        when "0101000001" => n11 <= "010001101100100101100101010101101010";
        when "0101000010" => n11 <= "010001100111010101100101010010001100";
        when "0101000011" => n11 <= "010001100010000101100101001110110000";
        when "0101000100" => n11 <= "010001011100110100100101001011010100";
        when "0101000101" => n11 <= "010001010111100011100101000111111001";
        when "0101000110" => n11 <= "010001010010010001100101000100011111";
        when "0101000111" => n11 <= "010001001100111110100101000001000111";
        when "0101001000" => n11 <= "010001000111101011100100111101101111";
        when "0101001001" => n11 <= "010001000010010111100100111010011000";
        when "0101001010" => n11 <= "010000111101000010100100110111000011";
        when "0101001011" => n11 <= "010000110111101101100100110011101110";
        when "0101001100" => n11 <= "010000110010010111100100110000011011";
        when "0101001101" => n11 <= "010000101101000000100100101101001000";
        when "0101001110" => n11 <= "010000100111101001100100101001110111";
        when "0101001111" => n11 <= "010000100010010001100100100110100111";
        when "0101010000" => n11 <= "010000011100111000100100100011010111";
        when "0101010001" => n11 <= "010000010111011111100100100000001001";
        when "0101010010" => n11 <= "010000010010000101100100011100111100";
        when "0101010011" => n11 <= "010000001100101010100100011001110000";
        when "0101010100" => n11 <= "010000000111001111100100010110100101";
        when "0101010101" => n11 <= "010000000001110100100100010011011011";
        when "0101010110" => n11 <= "001111111100010111100100010000010010";
        when "0101010111" => n11 <= "001111110110111010100100001101001010";
        when "0101011000" => n11 <= "001111110001011101100100001010000011";
        when "0101011001" => n11 <= "001111101011111110100100000110111110";
        when "0101011010" => n11 <= "001111100110100000100100000011111001";
        when "0101011011" => n11 <= "001111100001000000100100000000110110";
        when "0101011100" => n11 <= "001111011011100000100011111101110011";
        when "0101011101" => n11 <= "001111010110000000100011111010110010";
        when "0101011110" => n11 <= "001111010000011111100011110111110010";
        when "0101011111" => n11 <= "001111001010111101100011110100110010";
        when "0101100000" => n11 <= "001111000101011010100011110001110100";
        when "0101100001" => n11 <= "001110111111110111100011101110110111";
        when "0101100010" => n11 <= "001110111010010100100011101011111011";
        when "0101100011" => n11 <= "001110110100110000100011101001000001";
        when "0101100100" => n11 <= "001110101111001011100011100110000111";
        when "0101100101" => n11 <= "001110101001100110100011100011001110";
        when "0101100110" => n11 <= "001110100100000000100011100000010111";
        when "0101100111" => n11 <= "001110011110011010100011011101100000";
        when "0101101000" => n11 <= "001110011000110011100011011010101011";
        when "0101101001" => n11 <= "001110010011001011100011010111110111";
        when "0101101010" => n11 <= "001110001101100011100011010101000011";
        when "0101101011" => n11 <= "001110000111111011100011010010010001";
        when "0101101100" => n11 <= "001110000010010010100011001111100000";
        when "0101101101" => n11 <= "001101111100101000100011001100110001";
        when "0101101110" => n11 <= "001101110110111110100011001010000010";
        when "0101101111" => n11 <= "001101110001010011100011000111010100";
        when "0101110000" => n11 <= "001101101011101000100011000100101000";
        when "0101110001" => n11 <= "001101100101111100100011000001111100";
        when "0101110010" => n11 <= "001101100000010000100010111111010010";
        when "0101110011" => n11 <= "001101011010100011100010111100101001";
        when "0101110100" => n11 <= "001101010100110110100010111010000001";
        when "0101110101" => n11 <= "001101001111001000100010110111011010";
        when "0101110110" => n11 <= "001101001001011010100010110100110100";
        when "0101110111" => n11 <= "001101000011101011100010110010010000";
        when "0101111000" => n11 <= "001100111101111011100010101111101100";
        when "0101111001" => n11 <= "001100111000001011100010101101001010";
        when "0101111010" => n11 <= "001100110010011011100010101010101001";
        when "0101111011" => n11 <= "001100101100101010100010101000001000";
        when "0101111100" => n11 <= "001100100110111001100010100101101001";
        when "0101111101" => n11 <= "001100100001000111100010100011001100";
        when "0101111110" => n11 <= "001100011011010101100010100000101111";
        when "0101111111" => n11 <= "001100010101100010100010011110010011";
        when "0110000000" => n11 <= "001100001111101111100010011011111001";
        when "0110000001" => n11 <= "001100001001111011100010011001011111";
        when "0110000010" => n11 <= "001100000100000111100010010111000111";
        when "0110000011" => n11 <= "001011111110010010100010010100110000";
        when "0110000100" => n11 <= "001011111000011101100010010010011010";
        when "0110000101" => n11 <= "001011110010100111100010010000000110";
        when "0110000110" => n11 <= "001011101100110001100010001101110010";
        when "0110000111" => n11 <= "001011100110111011100010001011100000";
        when "0110001000" => n11 <= "001011100001000100100010001001001110";
        when "0110001001" => n11 <= "001011011011001100100010000110111110";
        when "0110001010" => n11 <= "001011010101010100100010000100101111";
        when "0110001011" => n11 <= "001011001111011100100010000010100001";
        when "0110001100" => n11 <= "001011001001100011100010000000010101";
        when "0110001101" => n11 <= "001011000011101010100001111110001001";
        when "0110001110" => n11 <= "001010111101110001100001111011111111";
        when "0110001111" => n11 <= "001010110111110111100001111001110101";
        when "0110010000" => n11 <= "001010110001111100100001110111101101";
        when "0110010001" => n11 <= "001010101100000010100001110101100111";
        when "0110010010" => n11 <= "001010100110000110100001110011100001";
        when "0110010011" => n11 <= "001010100000001011100001110001011100";
        when "0110010100" => n11 <= "001010011010001111100001101111011001";
        when "0110010101" => n11 <= "001010010100010010100001101101010111";
        when "0110010110" => n11 <= "001010001110010101100001101011010110";
        when "0110010111" => n11 <= "001010001000011000100001101001010110";
        when "0110011000" => n11 <= "001010000010011010100001100111010111";
        when "0110011001" => n11 <= "001001111100011100100001100101011001";
        when "0110011010" => n11 <= "001001110110011110100001100011011101";
        when "0110011011" => n11 <= "001001110000011111100001100001100010";
        when "0110011100" => n11 <= "001001101010100000100001011111101000";
        when "0110011101" => n11 <= "001001100100100000100001011101101111";
        when "0110011110" => n11 <= "001001011110100001100001011011110111";
        when "0110011111" => n11 <= "001001011000100000100001011010000001";
        when "0110100000" => n11 <= "001001010010100000100001011000001011";
        when "0110100001" => n11 <= "001001001100011111100001010110010111";
        when "0110100010" => n11 <= "001001000110011101100001010100100100";
        when "0110100011" => n11 <= "001001000000011100100001010010110011";
        when "0110100100" => n11 <= "001000111010011010100001010001000010";
        when "0110100101" => n11 <= "001000110100010111100001001111010011";
        when "0110100110" => n11 <= "001000101110010101100001001101100100";
        when "0110100111" => n11 <= "001000101000010001100001001011110111";
        when "0110101000" => n11 <= "001000100010001110100001001010001011";
        when "0110101001" => n11 <= "001000011100001010100001001000100001";
        when "0110101010" => n11 <= "001000010110000110100001000110110111";
        when "0110101011" => n11 <= "001000010000000010100001000101001111";
        when "0110101100" => n11 <= "001000001001111101100001000011101000";
        when "0110101101" => n11 <= "001000000011111000100001000010000010";
        when "0110101110" => n11 <= "000111111101110011100001000000011101";
        when "0110101111" => n11 <= "000111110111101101100000111110111010";
        when "0110110000" => n11 <= "000111110001100111100000111101011000";
        when "0110110001" => n11 <= "000111101011100001100000111011110110";
        when "0110110010" => n11 <= "000111100101011011100000111010010111";
        when "0110110011" => n11 <= "000111011111010100100000111000111000";
        when "0110110100" => n11 <= "000111011001001101100000110111011010";
        when "0110110101" => n11 <= "000111010011000101100000110101111110";
        when "0110110110" => n11 <= "000111001100111110100000110100100011";
        when "0110110111" => n11 <= "000111000110110110100000110011001001";
        when "0110111000" => n11 <= "000111000000101110100000110001110000";
        when "0110111001" => n11 <= "000110111010100101100000110000011001";
        when "0110111010" => n11 <= "000110110100011100100000101111000010";
        when "0110111011" => n11 <= "000110101110010011100000101101101101";
        when "0110111100" => n11 <= "000110101000001010100000101100011001";
        when "0110111101" => n11 <= "000110100010000000100000101011000111";
        when "0110111110" => n11 <= "000110011011110111100000101001110101";
        when "0110111111" => n11 <= "000110010101101101100000101000100101";
        when "0111000000" => n11 <= "000110001111100010100000100111010110";
        when "0111000001" => n11 <= "000110001001011000100000100110001000";
        when "0111000010" => n11 <= "000110000011001101100000100100111100";
        when "0111000011" => n11 <= "000101111101000010100000100011110000";
        when "0111000100" => n11 <= "000101110110110111100000100010100110";
        when "0111000101" => n11 <= "000101110000101011100000100001011101";
        when "0111000110" => n11 <= "000101101010100000100000100000010101";
        when "0111000111" => n11 <= "000101100100010100100000011111001111";
        when "0111001000" => n11 <= "000101011110001000100000011110001001";
        when "0111001001" => n11 <= "000101010111111100100000011101000101";
        when "0111001010" => n11 <= "000101010001101111100000011100000010";
        when "0111001011" => n11 <= "000101001011100010100000011011000000";
        when "0111001100" => n11 <= "000101000101010101100000011010000000";
        when "0111001101" => n11 <= "000100111111001000100000011001000001";
        when "0111001110" => n11 <= "000100111000111011100000011000000011";
        when "0111001111" => n11 <= "000100110010101101100000010111000110";
        when "0111010000" => n11 <= "000100101100100000100000010110001010";
        when "0111010001" => n11 <= "000100100110010010100000010101010000";
        when "0111010010" => n11 <= "000100100000000100100000010100010111";
        when "0111010011" => n11 <= "000100011001110110100000010011011111";
        when "0111010100" => n11 <= "000100010011100111100000010010101000";
        when "0111010101" => n11 <= "000100001101011001100000010001110010";
        when "0111010110" => n11 <= "000100000111001010100000010000111110";
        when "0111010111" => n11 <= "000100000000111011100000010000001011";
        when "0111011000" => n11 <= "000011111010101100100000001111011001";
        when "0111011001" => n11 <= "000011110100011101100000001110101001";
        when "0111011010" => n11 <= "000011101110001110100000001101111001";
        when "0111011011" => n11 <= "000011100111111110100000001101001011";
        when "0111011100" => n11 <= "000011100001101111100000001100011110";
        when "0111011101" => n11 <= "000011011011011111100000001011110010";
        when "0111011110" => n11 <= "000011010101001111100000001011001000";
        when "0111011111" => n11 <= "000011001110111111100000001010011111";
        when "0111100000" => n11 <= "000011001000101111100000001001110111";
        when "0111100001" => n11 <= "000011000010011111100000001001010000";
        when "0111100010" => n11 <= "000010111100001110100000001000101010";
        when "0111100011" => n11 <= "000010110101111110100000001000000110";
        when "0111100100" => n11 <= "000010101111101101100000000111100011";
        when "0111100101" => n11 <= "000010101001011100100000000111000001";
        when "0111100110" => n11 <= "000010100011001100100000000110100000";
        when "0111100111" => n11 <= "000010011100111011100000000110000001";
        when "0111101000" => n11 <= "000010010110101010100000000101100011";
        when "0111101001" => n11 <= "000010010000011001100000000101000110";
        when "0111101010" => n11 <= "000010001010001000100000000100101010";
        when "0111101011" => n11 <= "000010000011110110100000000100001111";
        when "0111101100" => n11 <= "000001111101100101100000000011110110";
        when "0111101101" => n11 <= "000001110111010100100000000011011110";
        when "0111101110" => n11 <= "000001110001000010100000000011000111";
        when "0111101111" => n11 <= "000001101010110001100000000010110010";
        when "0111110000" => n11 <= "000001100100011111100000000010011101";
        when "0111110001" => n11 <= "000001011110001101100000000010001010";
        when "0111110010" => n11 <= "000001010111111100100000000001111000";
        when "0111110011" => n11 <= "000001010001101010100000000001101000";
        when "0111110100" => n11 <= "000001001011011000100000000001011000";
        when "0111110101" => n11 <= "000001000101000110100000000001001010";
        when "0111110110" => n11 <= "000000111110110100100000000000111101";
        when "0111110111" => n11 <= "000000111000100010100000000000110001";
        when "0111111000" => n11 <= "000000110010010000100000000000100111";
        when "0111111001" => n11 <= "000000101011111110100000000000011110";
        when "0111111010" => n11 <= "000000100101101100100000000000010110";
        when "0111111011" => n11 <= "000000011111011010100000000000001111";
        when "0111111100" => n11 <= "000000011001001000100000000000001001";
        when "0111111101" => n11 <= "000000010010110110100000000000000101";
        when "0111111110" => n11 <= "000000001100100100100000000000000010";
        when "0111111111" => n11 <= "000000000110010010100000000000000000";
        when "1000000000" => n11 <= "000000000000000000100000000000000000";
        when "1000000001" => n11 <= "111111111001101101100000000000000000";
        when "1000000010" => n11 <= "111111110011011011100000000000000010";
        when "1000000011" => n11 <= "111111101101001001100000000000000101";
        when "1000000100" => n11 <= "111111100110110111100000000000001001";
        when "1000000101" => n11 <= "111111100000100101100000000000001111";
        when "1000000110" => n11 <= "111111011010010011100000000000010110";
        when "1000000111" => n11 <= "111111010100000001100000000000011110";
        when "1000001000" => n11 <= "111111001101101111100000000000100111";
        when "1000001001" => n11 <= "111111000111011101100000000000110001";
        when "1000001010" => n11 <= "111111000001001011100000000000111101";
        when "1000001011" => n11 <= "111110111010111001100000000001001010";
        when "1000001100" => n11 <= "111110110100100111100000000001011000";
        when "1000001101" => n11 <= "111110101110010101100000000001101000";
        when "1000001110" => n11 <= "111110101000000011100000000001111000";
        when "1000001111" => n11 <= "111110100001110010100000000010001010";
        when "1000010000" => n11 <= "111110011011100000100000000010011101";
        when "1000010001" => n11 <= "111110010101001110100000000010110010";
        when "1000010010" => n11 <= "111110001110111101100000000011000111";
        when "1000010011" => n11 <= "111110001000101011100000000011011110";
        when "1000010100" => n11 <= "111110000010011010100000000011110110";
        when "1000010101" => n11 <= "111101111100001001100000000100001111";
        when "1000010110" => n11 <= "111101110101110111100000000100101010";
        when "1000010111" => n11 <= "111101101111100110100000000101000110";
        when "1000011000" => n11 <= "111101101001010101100000000101100011";
        when "1000011001" => n11 <= "111101100011000100100000000110000001";
        when "1000011010" => n11 <= "111101011100110011100000000110100000";
        when "1000011011" => n11 <= "111101010110100011100000000111000001";
        when "1000011100" => n11 <= "111101010000010010100000000111100011";
        when "1000011101" => n11 <= "111101001010000001100000001000000110";
        when "1000011110" => n11 <= "111101000011110001100000001000101010";
        when "1000011111" => n11 <= "111100111101100000100000001001010000";
        when "1000100000" => n11 <= "111100110111010000100000001001110111";
        when "1000100001" => n11 <= "111100110001000000100000001010011111";
        when "1000100010" => n11 <= "111100101010110000100000001011001000";
        when "1000100011" => n11 <= "111100100100100000100000001011110010";
        when "1000100100" => n11 <= "111100011110010000100000001100011110";
        when "1000100101" => n11 <= "111100011000000001100000001101001011";
        when "1000100110" => n11 <= "111100010001110001100000001101111001";
        when "1000100111" => n11 <= "111100001011100010100000001110101001";
        when "1000101000" => n11 <= "111100000101010011100000001111011001";
        when "1000101001" => n11 <= "111011111111000100100000010000001011";
        when "1000101010" => n11 <= "111011111000110101100000010000111110";
        when "1000101011" => n11 <= "111011110010100110100000010001110010";
        when "1000101100" => n11 <= "111011101100011000100000010010101000";
        when "1000101101" => n11 <= "111011100110001001100000010011011111";
        when "1000101110" => n11 <= "111011011111111011100000010100010111";
        when "1000101111" => n11 <= "111011011001101101100000010101010000";
        when "1000110000" => n11 <= "111011010011011111100000010110001010";
        when "1000110001" => n11 <= "111011001101010010100000010111000110";
        when "1000110010" => n11 <= "111011000111000100100000011000000011";
        when "1000110011" => n11 <= "111011000000110111100000011001000001";
        when "1000110100" => n11 <= "111010111010101010100000011010000000";
        when "1000110101" => n11 <= "111010110100011101100000011011000000";
        when "1000110110" => n11 <= "111010101110010000100000011100000010";
        when "1000110111" => n11 <= "111010101000000011100000011101000101";
        when "1000111000" => n11 <= "111010100001110111100000011110001001";
        when "1000111001" => n11 <= "111010011011101011100000011111001111";
        when "1000111010" => n11 <= "111010010101011111100000100000010101";
        when "1000111011" => n11 <= "111010001111010100100000100001011101";
        when "1000111100" => n11 <= "111010001001001000100000100010100110";
        when "1000111101" => n11 <= "111010000010111101100000100011110000";
        when "1000111110" => n11 <= "111001111100110010100000100100111100";
        when "1000111111" => n11 <= "111001110110100111100000100110001000";
        when "1001000000" => n11 <= "111001110000011101100000100111010110";
        when "1001000001" => n11 <= "111001101010010010100000101000100101";
        when "1001000010" => n11 <= "111001100100001000100000101001110101";
        when "1001000011" => n11 <= "111001011101111111100000101011000111";
        when "1001000100" => n11 <= "111001010111110101100000101100011001";
        when "1001000101" => n11 <= "111001010001101100100000101101101101";
        when "1001000110" => n11 <= "111001001011100011100000101111000010";
        when "1001000111" => n11 <= "111001000101011010100000110000011001";
        when "1001001000" => n11 <= "111000111111010001100000110001110000";
        when "1001001001" => n11 <= "111000111001001001100000110011001001";
        when "1001001010" => n11 <= "111000110011000001100000110100100011";
        when "1001001011" => n11 <= "111000101100111010100000110101111110";
        when "1001001100" => n11 <= "111000100110110010100000110111011010";
        when "1001001101" => n11 <= "111000100000101011100000111000111000";
        when "1001001110" => n11 <= "111000011010100100100000111010010111";
        when "1001001111" => n11 <= "111000010100011110100000111011110110";
        when "1001010000" => n11 <= "111000001110011000100000111101011000";
        when "1001010001" => n11 <= "111000001000010010100000111110111010";
        when "1001010010" => n11 <= "111000000010001100100001000000011101";
        when "1001010011" => n11 <= "110111111100000111100001000010000010";
        when "1001010100" => n11 <= "110111110110000010100001000011101000";
        when "1001010101" => n11 <= "110111101111111101100001000101001111";
        when "1001010110" => n11 <= "110111101001111001100001000110110111";
        when "1001010111" => n11 <= "110111100011110101100001001000100001";
        when "1001011000" => n11 <= "110111011101110001100001001010001011";
        when "1001011001" => n11 <= "110111010111101110100001001011110111";
        when "1001011010" => n11 <= "110111010001101010100001001101100100";
        when "1001011011" => n11 <= "110111001011101000100001001111010011";
        when "1001011100" => n11 <= "110111000101100101100001010001000010";
        when "1001011101" => n11 <= "110110111111100011100001010010110011";
        when "1001011110" => n11 <= "110110111001100010100001010100100100";
        when "1001011111" => n11 <= "110110110011100000100001010110010111";
        when "1001100000" => n11 <= "110110101101011111100001011000001011";
        when "1001100001" => n11 <= "110110100111011111100001011010000001";
        when "1001100010" => n11 <= "110110100001011110100001011011110111";
        when "1001100011" => n11 <= "110110011011011111100001011101101111";
        when "1001100100" => n11 <= "110110010101011111100001011111101000";
        when "1001100101" => n11 <= "110110001111100000100001100001100010";
        when "1001100110" => n11 <= "110110001001100001100001100011011101";
        when "1001100111" => n11 <= "110110000011100011100001100101011001";
        when "1001101000" => n11 <= "110101111101100101100001100111010111";
        when "1001101001" => n11 <= "110101110111100111100001101001010110";
        when "1001101010" => n11 <= "110101110001101010100001101011010110";
        when "1001101011" => n11 <= "110101101011101101100001101101010111";
        when "1001101100" => n11 <= "110101100101110000100001101111011001";
        when "1001101101" => n11 <= "110101011111110100100001110001011100";
        when "1001101110" => n11 <= "110101011001111001100001110011100001";
        when "1001101111" => n11 <= "110101010011111101100001110101100111";
        when "1001110000" => n11 <= "110101001110000011100001110111101101";
        when "1001110001" => n11 <= "110101001000001000100001111001110101";
        when "1001110010" => n11 <= "110101000010001110100001111011111111";
        when "1001110011" => n11 <= "110100111100010101100001111110001001";
        when "1001110100" => n11 <= "110100110110011100100010000000010101";
        when "1001110101" => n11 <= "110100110000100011100010000010100001";
        when "1001110110" => n11 <= "110100101010101011100010000100101111";
        when "1001110111" => n11 <= "110100100100110011100010000110111110";
        when "1001111000" => n11 <= "110100011110111011100010001001001110";
        when "1001111001" => n11 <= "110100011001000100100010001011100000";
        when "1001111010" => n11 <= "110100010011001110100010001101110010";
        when "1001111011" => n11 <= "110100001101011000100010010000000110";
        when "1001111100" => n11 <= "110100000111100010100010010010011010";
        when "1001111101" => n11 <= "110100000001101101100010010100110000";
        when "1001111110" => n11 <= "110011111011111000100010010111000111";
        when "1001111111" => n11 <= "110011110110000100100010011001011111";
        when "1010000000" => n11 <= "110011110000010000100010011011111001";
        when "1010000001" => n11 <= "110011101010011101100010011110010011";
        when "1010000010" => n11 <= "110011100100101010100010100000101111";
        when "1010000011" => n11 <= "110011011110111000100010100011001100";
        when "1010000100" => n11 <= "110011011001000110100010100101101001";
        when "1010000101" => n11 <= "110011010011010101100010101000001000";
        when "1010000110" => n11 <= "110011001101100100100010101010101001";
        when "1010000111" => n11 <= "110011000111110100100010101101001010";
        when "1010001000" => n11 <= "110011000010000100100010101111101100";
        when "1010001001" => n11 <= "110010111100010100100010110010010000";
        when "1010001010" => n11 <= "110010110110100101100010110100110100";
        when "1010001011" => n11 <= "110010110000110111100010110111011010";
        when "1010001100" => n11 <= "110010101011001001100010111010000001";
        when "1010001101" => n11 <= "110010100101011100100010111100101001";
        when "1010001110" => n11 <= "110010011111101111100010111111010010";
        when "1010001111" => n11 <= "110010011010000011100011000001111100";
        when "1010010000" => n11 <= "110010010100010111100011000100101000";
        when "1010010001" => n11 <= "110010001110101100100011000111010100";
        when "1010010010" => n11 <= "110010001001000001100011001010000010";
        when "1010010011" => n11 <= "110010000011010111100011001100110001";
        when "1010010100" => n11 <= "110001111101101101100011001111100000";
        when "1010010101" => n11 <= "110001111000000100100011010010010001";
        when "1010010110" => n11 <= "110001110010011100100011010101000011";
        when "1010010111" => n11 <= "110001101100110100100011010111110111";
        when "1010011000" => n11 <= "110001100111001100100011011010101011";
        when "1010011001" => n11 <= "110001100001100101100011011101100000";
        when "1010011010" => n11 <= "110001011011111111100011100000010111";
        when "1010011011" => n11 <= "110001010110011001100011100011001110";
        when "1010011100" => n11 <= "110001010000110100100011100110000111";
        when "1010011101" => n11 <= "110001001011001111100011101001000001";
        when "1010011110" => n11 <= "110001000101101011100011101011111011";
        when "1010011111" => n11 <= "110001000000001000100011101110110111";
        when "1010100000" => n11 <= "110000111010100101100011110001110100";
        when "1010100001" => n11 <= "110000110101000010100011110100110010";
        when "1010100010" => n11 <= "110000101111100000100011110111110010";
        when "1010100011" => n11 <= "110000101001111111100011111010110010";
        when "1010100100" => n11 <= "110000100100011111100011111101110011";
        when "1010100101" => n11 <= "110000011110111111100100000000110110";
        when "1010100110" => n11 <= "110000011001011111100100000011111001";
        when "1010100111" => n11 <= "110000010100000001100100000110111110";
        when "1010101000" => n11 <= "110000001110100010100100001010000011";
        when "1010101001" => n11 <= "110000001001000101100100001101001010";
        when "1010101010" => n11 <= "110000000011101000100100010000010010";
        when "1010101011" => n11 <= "101111111110001011100100010011011011";
        when "1010101100" => n11 <= "101111111000110000100100010110100101";
        when "1010101101" => n11 <= "101111110011010101100100011001110000";
        when "1010101110" => n11 <= "101111101101111010100100011100111100";
        when "1010101111" => n11 <= "101111101000100000100100100000001001";
        when "1010110000" => n11 <= "101111100011000111100100100011010111";
        when "1010110001" => n11 <= "101111011101101110100100100110100111";
        when "1010110010" => n11 <= "101111011000010110100100101001110111";
        when "1010110011" => n11 <= "101111010010111111100100101101001000";
        when "1010110100" => n11 <= "101111001101101000100100110000011011";
        when "1010110101" => n11 <= "101111001000010010100100110011101110";
        when "1010110110" => n11 <= "101111000010111101100100110111000011";
        when "1010110111" => n11 <= "101110111101101000100100111010011000";
        when "1010111000" => n11 <= "101110111000010100100100111101101111";
        when "1010111001" => n11 <= "101110110011000001100101000001000111";
        when "1010111010" => n11 <= "101110101101101110100101000100011111";
        when "1010111011" => n11 <= "101110101000011100100101000111111001";
        when "1010111100" => n11 <= "101110100011001011100101001011010100";
        when "1010111101" => n11 <= "101110011101111010100101001110110000";
        when "1010111110" => n11 <= "101110011000101010100101010010001100";
        when "1010111111" => n11 <= "101110010011011010100101010101101010";
        when "1011000000" => n11 <= "101110001110001100100101011001001001";
        when "1011000001" => n11 <= "101110001000111110100101011100101001";
        when "1011000010" => n11 <= "101110000011110000100101100000001010";
        when "1011000011" => n11 <= "101101111110100100100101100011101100";
        when "1011000100" => n11 <= "101101111001011000100101100111001111";
        when "1011000101" => n11 <= "101101110100001101100101101010110011";
        when "1011000110" => n11 <= "101101101111000010100101101110011000";
        when "1011000111" => n11 <= "101101101001111000100101110001111110";
        when "1011001000" => n11 <= "101101100100101111100101110101100101";
        when "1011001001" => n11 <= "101101011111100111100101111001001101";
        when "1011001010" => n11 <= "101101011010011111100101111100110110";
        when "1011001011" => n11 <= "101101010101011000100110000000100000";
        when "1011001100" => n11 <= "101101010000010010100110000100001011";
        when "1011001101" => n11 <= "101101001011001100100110000111110111";
        when "1011001110" => n11 <= "101101000110000111100110001011100100";
        when "1011001111" => n11 <= "101101000001000011100110001111010010";
        when "1011010000" => n11 <= "101100111100000000100110010011000001";
        when "1011010001" => n11 <= "101100110110111101100110010110110010";
        when "1011010010" => n11 <= "101100110001111011100110011010100011";
        when "1011010011" => n11 <= "101100101100111010100110011110010101";
        when "1011010100" => n11 <= "101100100111111010100110100010001000";
        when "1011010101" => n11 <= "101100100010111010100110100101111100";
        when "1011010110" => n11 <= "101100011101111011100110101001110001";
        when "1011010111" => n11 <= "101100011000111101100110101101100110";
        when "1011011000" => n11 <= "101100010100000000100110110001011101";
        when "1011011001" => n11 <= "101100001111000011100110110101010101";
        when "1011011010" => n11 <= "101100001010000111100110111001001110";
        when "1011011011" => n11 <= "101100000101001100100110111101001000";
        when "1011011100" => n11 <= "101100000000010010100111000001000011";
        when "1011011101" => n11 <= "101011111011011000100111000100111110";
        when "1011011110" => n11 <= "101011110110100000100111001000111011";
        when "1011011111" => n11 <= "101011110001101000100111001100111001";
        when "1011100000" => n11 <= "101011101100110000100111010000110111";
        when "1011100001" => n11 <= "101011100111111010100111010100110111";
        when "1011100010" => n11 <= "101011100011000100100111011000111000";
        when "1011100011" => n11 <= "101011011110001111100111011100111001";
        when "1011100100" => n11 <= "101011011001011011100111100000111011";
        when "1011100101" => n11 <= "101011010100101000100111100100111111";
        when "1011100110" => n11 <= "101011001111110101100111101001000011";
        when "1011100111" => n11 <= "101011001011000100100111101101001000";
        when "1011101000" => n11 <= "101011000110010011100111110001001111";
        when "1011101001" => n11 <= "101011000001100011100111110101010110";
        when "1011101010" => n11 <= "101010111100110011100111111001011110";
        when "1011101011" => n11 <= "101010111000000101100111111101100111";
        when "1011101100" => n11 <= "101010110011010111101000000001110001";
        when "1011101101" => n11 <= "101010101110101011101000000101111100";
        when "1011101110" => n11 <= "101010101001111110101000001010000111";
        when "1011101111" => n11 <= "101010100101010011101000001110010100";
        when "1011110000" => n11 <= "101010100000101001101000010010100010";
        when "1011110001" => n11 <= "101010011011111111101000010110110000";
        when "1011110010" => n11 <= "101010010111010111101000011010111111";
        when "1011110011" => n11 <= "101010010010101111101000011111010000";
        when "1011110100" => n11 <= "101010001110001000101000100011100001";
        when "1011110101" => n11 <= "101010001001100010101000100111110011";
        when "1011110110" => n11 <= "101010000100111100101000101100000110";
        when "1011110111" => n11 <= "101010000000011000101000110000011010";
        when "1011111000" => n11 <= "101001111011110100101000110100101111";
        when "1011111001" => n11 <= "101001110111010001101000111001000101";
        when "1011111010" => n11 <= "101001110010101111101000111101011011";
        when "1011111011" => n11 <= "101001101110001110101001000001110011";
        when "1011111100" => n11 <= "101001101001101110101001000110001011";
        when "1011111101" => n11 <= "101001100101001111101001001010100101";
        when "1011111110" => n11 <= "101001100000110000101001001110111111";
        when "1011111111" => n11 <= "101001011100010010101001010011011010";
        when "1100000000" => n11 <= "101001010111110110101001010111110110";
        when "1100000001" => n11 <= "101001010011011010101001011100010010";
        when "1100000010" => n11 <= "101001001110111111101001100000110000";
        when "1100000011" => n11 <= "101001001010100101101001100101001111";
        when "1100000100" => n11 <= "101001000110001011101001101001101110";
        when "1100000101" => n11 <= "101001000001110011101001101110001110";
        when "1100000110" => n11 <= "101000111101011011101001110010101111";
        when "1100000111" => n11 <= "101000111001000101101001110111010001";
        when "1100001000" => n11 <= "101000110100101111101001111011110100";
        when "1100001001" => n11 <= "101000110000011010101010000000011000";
        when "1100001010" => n11 <= "101000101100000110101010000100111100";
        when "1100001011" => n11 <= "101000100111110011101010001001100010";
        when "1100001100" => n11 <= "101000100011100001101010001110001000";
        when "1100001101" => n11 <= "101000011111010000101010010010101111";
        when "1100001110" => n11 <= "101000011010111111101010010111010111";
        when "1100001111" => n11 <= "101000010110110000101010011011111111";
        when "1100010000" => n11 <= "101000010010100010101010100000101001";
        when "1100010001" => n11 <= "101000001110010100101010100101010011";
        when "1100010010" => n11 <= "101000001010000111101010101001111110";
        when "1100010011" => n11 <= "101000000101111100101010101110101011";
        when "1100010100" => n11 <= "101000000001110001101010110011010111";
        when "1100010101" => n11 <= "100111111101100111101010111000000101";
        when "1100010110" => n11 <= "100111111001011110101010111100110011";
        when "1100010111" => n11 <= "100111110101010110101011000001100011";
        when "1100011000" => n11 <= "100111110001001111101011000110010011";
        when "1100011001" => n11 <= "100111101101001000101011001011000100";
        when "1100011010" => n11 <= "100111101001000011101011001111110101";
        when "1100011011" => n11 <= "100111100100111111101011010100101000";
        when "1100011100" => n11 <= "100111100000111011101011011001011011";
        when "1100011101" => n11 <= "100111011100111001101011011110001111";
        when "1100011110" => n11 <= "100111011000111000101011100011000100";
        when "1100011111" => n11 <= "100111010100110111101011100111111010";
        when "1100100000" => n11 <= "100111010000110111101011101100110000";
        when "1100100001" => n11 <= "100111001100111001101011110001101000";
        when "1100100010" => n11 <= "100111001000111011101011110110100000";
        when "1100100011" => n11 <= "100111000100111110101011111011011000";
        when "1100100100" => n11 <= "100111000001000011101100000000010010";
        when "1100100101" => n11 <= "100110111101001000101100000101001100";
        when "1100100110" => n11 <= "100110111001001110101100001010000111";
        when "1100100111" => n11 <= "100110110101010101101100001111000011";
        when "1100101000" => n11 <= "100110110001011101101100010100000000";
        when "1100101001" => n11 <= "100110101101100110101100011000111101";
        when "1100101010" => n11 <= "100110101001110001101100011101111011";
        when "1100101011" => n11 <= "100110100101111100101100100010111010";
        when "1100101100" => n11 <= "100110100010001000101100100111111010";
        when "1100101101" => n11 <= "100110011110010101101100101100111010";
        when "1100101110" => n11 <= "100110011010100011101100110001111011";
        when "1100101111" => n11 <= "100110010110110010101100110110111101";
        when "1100110000" => n11 <= "100110010011000001101100111100000000";
        when "1100110001" => n11 <= "100110001111010010101101000001000011";
        when "1100110010" => n11 <= "100110001011100100101101000110000111";
        when "1100110011" => n11 <= "100110000111110111101101001011001100";
        when "1100110100" => n11 <= "100110000100001011101101010000010010";
        when "1100110101" => n11 <= "100110000000100000101101010101011000";
        when "1100110110" => n11 <= "100101111100110110101101011010011111";
        when "1100110111" => n11 <= "100101111001001101101101011111100111";
        when "1100111000" => n11 <= "100101110101100101101101100100101111";
        when "1100111001" => n11 <= "100101110001111110101101101001111000";
        when "1100111010" => n11 <= "100101101110011000101101101111000010";
        when "1100111011" => n11 <= "100101101010110011101101110100001101";
        when "1100111100" => n11 <= "100101100111001111101101111001011000";
        when "1100111101" => n11 <= "100101100011101100101101111110100100";
        when "1100111110" => n11 <= "100101100000001010101110000011110000";
        when "1100111111" => n11 <= "100101011100101001101110001000111110";
        when "1101000000" => n11 <= "100101011001001001101110001110001100";
        when "1101000001" => n11 <= "100101010101101010101110010011011010";
        when "1101000010" => n11 <= "100101010010001100101110011000101010";
        when "1101000011" => n11 <= "100101001110110000101110011101111010";
        when "1101000100" => n11 <= "100101001011010100101110100011001011";
        when "1101000101" => n11 <= "100101000111111001101110101000011100";
        when "1101000110" => n11 <= "100101000100011111101110101101101110";
        when "1101000111" => n11 <= "100101000001000111101110110011000001";
        when "1101001000" => n11 <= "100100111101101111101110111000010100";
        when "1101001001" => n11 <= "100100111010011000101110111101101000";
        when "1101001010" => n11 <= "100100110111000011101111000010111101";
        when "1101001011" => n11 <= "100100110011101110101111001000010010";
        when "1101001100" => n11 <= "100100110000011011101111001101101000";
        when "1101001101" => n11 <= "100100101101001000101111010010111111";
        when "1101001110" => n11 <= "100100101001110111101111011000010110";
        when "1101001111" => n11 <= "100100100110100111101111011101101110";
        when "1101010000" => n11 <= "100100100011010111101111100011000111";
        when "1101010001" => n11 <= "100100100000001001101111101000100000";
        when "1101010010" => n11 <= "100100011100111100101111101101111010";
        when "1101010011" => n11 <= "100100011001110000101111110011010101";
        when "1101010100" => n11 <= "100100010110100101101111111000110000";
        when "1101010101" => n11 <= "100100010011011011101111111110001011";
        when "1101010110" => n11 <= "100100010000010010110000000011101000";
        when "1101010111" => n11 <= "100100001101001010110000001001000101";
        when "1101011000" => n11 <= "100100001010000011110000001110100010";
        when "1101011001" => n11 <= "100100000110111110110000010100000001";
        when "1101011010" => n11 <= "100100000011111001110000011001011111";
        when "1101011011" => n11 <= "100100000000110110110000011110111111";
        when "1101011100" => n11 <= "100011111101110011110000100100011111";
        when "1101011101" => n11 <= "100011111010110010110000101001111111";
        when "1101011110" => n11 <= "100011110111110010110000101111100000";
        when "1101011111" => n11 <= "100011110100110010110000110101000010";
        when "1101100000" => n11 <= "100011110001110100110000111010100101";
        when "1101100001" => n11 <= "100011101110110111110001000000001000";
        when "1101100010" => n11 <= "100011101011111011110001000101101011";
        when "1101100011" => n11 <= "100011101001000001110001001011001111";
        when "1101100100" => n11 <= "100011100110000111110001010000110100";
        when "1101100101" => n11 <= "100011100011001110110001010110011001";
        when "1101100110" => n11 <= "100011100000010111110001011011111111";
        when "1101100111" => n11 <= "100011011101100000110001100001100101";
        when "1101101000" => n11 <= "100011011010101011110001100111001100";
        when "1101101001" => n11 <= "100011010111110111110001101100110100";
        when "1101101010" => n11 <= "100011010101000011110001110010011100";
        when "1101101011" => n11 <= "100011010010010001110001111000000100";
        when "1101101100" => n11 <= "100011001111100000110001111101101101";
        when "1101101101" => n11 <= "100011001100110001110010000011010111";
        when "1101101110" => n11 <= "100011001010000010110010001001000001";
        when "1101101111" => n11 <= "100011000111010100110010001110101100";
        when "1101110000" => n11 <= "100011000100101000110010010100010111";
        when "1101110001" => n11 <= "100011000001111100110010011010000011";
        when "1101110010" => n11 <= "100010111111010010110010011111101111";
        when "1101110011" => n11 <= "100010111100101001110010100101011100";
        when "1101110100" => n11 <= "100010111010000001110010101011001001";
        when "1101110101" => n11 <= "100010110111011010110010110000110111";
        when "1101110110" => n11 <= "100010110100110100110010110110100101";
        when "1101110111" => n11 <= "100010110010010000110010111100010100";
        when "1101111000" => n11 <= "100010101111101100110011000010000100";
        when "1101111001" => n11 <= "100010101101001010110011000111110100";
        when "1101111010" => n11 <= "100010101010101001110011001101100100";
        when "1101111011" => n11 <= "100010101000001000110011010011010101";
        when "1101111100" => n11 <= "100010100101101001110011011001000110";
        when "1101111101" => n11 <= "100010100011001100110011011110111000";
        when "1101111110" => n11 <= "100010100000101111110011100100101010";
        when "1101111111" => n11 <= "100010011110010011110011101010011101";
        when "1110000000" => n11 <= "100010011011111001110011110000010000";
        when "1110000001" => n11 <= "100010011001011111110011110110000100";
        when "1110000010" => n11 <= "100010010111000111110011111011111000";
        when "1110000011" => n11 <= "100010010100110000110100000001101101";
        when "1110000100" => n11 <= "100010010010011010110100000111100010";
        when "1110000101" => n11 <= "100010010000000110110100001101011000";
        when "1110000110" => n11 <= "100010001101110010110100010011001110";
        when "1110000111" => n11 <= "100010001011100000110100011001000100";
        when "1110001000" => n11 <= "100010001001001110110100011110111011";
        when "1110001001" => n11 <= "100010000110111110110100100100110011";
        when "1110001010" => n11 <= "100010000100101111110100101010101011";
        when "1110001011" => n11 <= "100010000010100001110100110000100011";
        when "1110001100" => n11 <= "100010000000010101110100110110011100";
        when "1110001101" => n11 <= "100001111110001001110100111100010101";
        when "1110001110" => n11 <= "100001111011111111110101000010001110";
        when "1110001111" => n11 <= "100001111001110101110101001000001000";
        when "1110010000" => n11 <= "100001110111101101110101001110000011";
        when "1110010001" => n11 <= "100001110101100111110101010011111101";
        when "1110010010" => n11 <= "100001110011100001110101011001111001";
        when "1110010011" => n11 <= "100001110001011100110101011111110100";
        when "1110010100" => n11 <= "100001101111011001110101100101110000";
        when "1110010101" => n11 <= "100001101101010111110101101011101101";
        when "1110010110" => n11 <= "100001101011010110110101110001101010";
        when "1110010111" => n11 <= "100001101001010110110101110111100111";
        when "1110011000" => n11 <= "100001100111010111110101111101100101";
        when "1110011001" => n11 <= "100001100101011001110110000011100011";
        when "1110011010" => n11 <= "100001100011011101110110001001100001";
        when "1110011011" => n11 <= "100001100001100010110110001111100000";
        when "1110011100" => n11 <= "100001011111101000110110010101011111";
        when "1110011101" => n11 <= "100001011101101111110110011011011111";
        when "1110011110" => n11 <= "100001011011110111110110100001011110";
        when "1110011111" => n11 <= "100001011010000001110110100111011111";
        when "1110100000" => n11 <= "100001011000001011110110101101011111";
        when "1110100001" => n11 <= "100001010110010111110110110011100000";
        when "1110100010" => n11 <= "100001010100100100110110111001100010";
        when "1110100011" => n11 <= "100001010010110011110110111111100011";
        when "1110100100" => n11 <= "100001010001000010110111000101100101";
        when "1110100101" => n11 <= "100001001111010011110111001011101000";
        when "1110100110" => n11 <= "100001001101100100110111010001101010";
        when "1110100111" => n11 <= "100001001011110111110111010111101110";
        when "1110101000" => n11 <= "100001001010001011110111011101110001";
        when "1110101001" => n11 <= "100001001000100001110111100011110101";
        when "1110101010" => n11 <= "100001000110110111110111101001111001";
        when "1110101011" => n11 <= "100001000101001111110111101111111101";
        when "1110101100" => n11 <= "100001000011101000110111110110000010";
        when "1110101101" => n11 <= "100001000010000010110111111100000111";
        when "1110101110" => n11 <= "100001000000011101111000000010001100";
        when "1110101111" => n11 <= "100000111110111010111000001000010010";
        when "1110110000" => n11 <= "100000111101011000111000001110011000";
        when "1110110001" => n11 <= "100000111011110110111000010100011110";
        when "1110110010" => n11 <= "100000111010010111111000011010100100";
        when "1110110011" => n11 <= "100000111000111000111000100000101011";
        when "1110110100" => n11 <= "100000110111011010111000100110110010";
        when "1110110101" => n11 <= "100000110101111110111000101100111010";
        when "1110110110" => n11 <= "100000110100100011111000110011000001";
        when "1110110111" => n11 <= "100000110011001001111000111001001001";
        when "1110111000" => n11 <= "100000110001110000111000111111010001";
        when "1110111001" => n11 <= "100000110000011001111001000101011010";
        when "1110111010" => n11 <= "100000101111000010111001001011100011";
        when "1110111011" => n11 <= "100000101101101101111001010001101100";
        when "1110111100" => n11 <= "100000101100011001111001010111110101";
        when "1110111101" => n11 <= "100000101011000111111001011101111111";
        when "1110111110" => n11 <= "100000101001110101111001100100001000";
        when "1110111111" => n11 <= "100000101000100101111001101010010010";
        when "1111000000" => n11 <= "100000100111010110111001110000011101";
        when "1111000001" => n11 <= "100000100110001000111001110110100111";
        when "1111000010" => n11 <= "100000100100111100111001111100110010";
        when "1111000011" => n11 <= "100000100011110000111010000010111101";
        when "1111000100" => n11 <= "100000100010100110111010001001001000";
        when "1111000101" => n11 <= "100000100001011101111010001111010100";
        when "1111000110" => n11 <= "100000100000010101111010010101011111";
        when "1111000111" => n11 <= "100000011111001111111010011011101011";
        when "1111001000" => n11 <= "100000011110001001111010100001110111";
        when "1111001001" => n11 <= "100000011101000101111010101000000011";
        when "1111001010" => n11 <= "100000011100000010111010101110010000";
        when "1111001011" => n11 <= "100000011011000000111010110100011101";
        when "1111001100" => n11 <= "100000011010000000111010111010101010";
        when "1111001101" => n11 <= "100000011001000001111011000000110111";
        when "1111001110" => n11 <= "100000011000000011111011000111000100";
        when "1111001111" => n11 <= "100000010111000110111011001101010010";
        when "1111010000" => n11 <= "100000010110001010111011010011011111";
        when "1111010001" => n11 <= "100000010101010000111011011001101101";
        when "1111010010" => n11 <= "100000010100010111111011011111111011";
        when "1111010011" => n11 <= "100000010011011111111011100110001001";
        when "1111010100" => n11 <= "100000010010101000111011101100011000";
        when "1111010101" => n11 <= "100000010001110010111011110010100110";
        when "1111010110" => n11 <= "100000010000111110111011111000110101";
        when "1111010111" => n11 <= "100000010000001011111011111111000100";
        when "1111011000" => n11 <= "100000001111011001111100000101010011";
        when "1111011001" => n11 <= "100000001110101001111100001011100010";
        when "1111011010" => n11 <= "100000001101111001111100010001110001";
        when "1111011011" => n11 <= "100000001101001011111100011000000001";
        when "1111011100" => n11 <= "100000001100011110111100011110010000";
        when "1111011101" => n11 <= "100000001011110010111100100100100000";
        when "1111011110" => n11 <= "100000001011001000111100101010110000";
        when "1111011111" => n11 <= "100000001010011111111100110001000000";
        when "1111100000" => n11 <= "100000001001110111111100110111010000";
        when "1111100001" => n11 <= "100000001001010000111100111101100000";
        when "1111100010" => n11 <= "100000001000101010111101000011110001";
        when "1111100011" => n11 <= "100000001000000110111101001010000001";
        when "1111100100" => n11 <= "100000000111100011111101010000010010";
        when "1111100101" => n11 <= "100000000111000001111101010110100011";
        when "1111100110" => n11 <= "100000000110100000111101011100110011";
        when "1111100111" => n11 <= "100000000110000001111101100011000100";
        when "1111101000" => n11 <= "100000000101100011111101101001010101";
        when "1111101001" => n11 <= "100000000101000110111101101111100110";
        when "1111101010" => n11 <= "100000000100101010111101110101110111";
        when "1111101011" => n11 <= "100000000100001111111101111100001001";
        when "1111101100" => n11 <= "100000000011110110111110000010011010";
        when "1111101101" => n11 <= "100000000011011110111110001000101011";
        when "1111101110" => n11 <= "100000000011000111111110001110111101";
        when "1111101111" => n11 <= "100000000010110010111110010101001110";
        when "1111110000" => n11 <= "100000000010011101111110011011100000";
        when "1111110001" => n11 <= "100000000010001010111110100001110010";
        when "1111110010" => n11 <= "100000000001111000111110101000000011";
        when "1111110011" => n11 <= "100000000001101000111110101110010101";
        when "1111110100" => n11 <= "100000000001011000111110110100100111";
        when "1111110101" => n11 <= "100000000001001010111110111010111001";
        when "1111110110" => n11 <= "100000000000111101111111000001001011";
        when "1111110111" => n11 <= "100000000000110001111111000111011101";
        when "1111111000" => n11 <= "100000000000100111111111001101101111";
        when "1111111001" => n11 <= "100000000000011110111111010100000001";
        when "1111111010" => n11 <= "100000000000010110111111011010010011";
        when "1111111011" => n11 <= "100000000000001111111111100000100101";
        when "1111111100" => n11 <= "100000000000001001111111100110110111";
        when "1111111101" => n11 <= "100000000000000101111111101101001001";
        when "1111111110" => n11 <= "100000000000000010111111110011011011";
        when "1111111111" => n11 <= "100000000000000000111111111001101101";
        when others => n11 <= "XXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX";
      end case;
    end if;
  end if;
end process;
n12 <= n11(35 downto 35) &
  n11(34 downto 34) &
  n11(33 downto 33) &
  n11(32 downto 32) &
  n11(31 downto 31) &
  n11(30 downto 30) &
  n11(29 downto 29) &
  n11(28 downto 28) &
  n11(27 downto 27) &
  n11(26 downto 26) &
  n11(25 downto 25) &
  n11(24 downto 24) &
  n11(23 downto 23) &
  n11(22 downto 22) &
  n11(21 downto 21) &
  n11(20 downto 20) &
  n11(19 downto 19) &
  n11(18 downto 18);
n13 <= n11(17 downto 17) &
  n11(16 downto 16) &
  n11(15 downto 15) &
  n11(14 downto 14) &
  n11(13 downto 13) &
  n11(12 downto 12) &
  n11(11 downto 11) &
  n11(10 downto 10) &
  n11(9 downto 9) &
  n11(8 downto 8) &
  n11(7 downto 7) &
  n11(6 downto 6) &
  n11(5 downto 5) &
  n11(4 downto 4) &
  n11(3 downto 3) &
  n11(2 downto 2) &
  n11(1 downto 1) &
  n11(0 downto 0);
n14 <= unsigned(signed(n5) * signed(n12));
n15 <= n14(34 downto 34) &
  n14(33 downto 33) &
  n14(32 downto 32) &
  n14(31 downto 31) &
  n14(30 downto 30) &
  n14(29 downto 29) &
  n14(28 downto 28) &
  n14(27 downto 27) &
  n14(26 downto 26) &
  n14(25 downto 25) &
  n14(24 downto 24) &
  n14(23 downto 23) &
  n14(22 downto 22) &
  n14(21 downto 21) &
  n14(20 downto 20) &
  n14(19 downto 19) &
  n14(18 downto 18) &
  n14(17 downto 17);
process (clock_c) begin
  if rising_edge(clock_c) then
    if i5 = "1" then
      n16 <= "000000000000000000";
    elsif i4 = "1" then
      n16 <= n15;
    end if;
  end if;
end process;
n17 <= unsigned(signed(n6) * signed(n13));
n18 <= n17(34 downto 34) &
  n17(33 downto 33) &
  n17(32 downto 32) &
  n17(31 downto 31) &
  n17(30 downto 30) &
  n17(29 downto 29) &
  n17(28 downto 28) &
  n17(27 downto 27) &
  n17(26 downto 26) &
  n17(25 downto 25) &
  n17(24 downto 24) &
  n17(23 downto 23) &
  n17(22 downto 22) &
  n17(21 downto 21) &
  n17(20 downto 20) &
  n17(19 downto 19) &
  n17(18 downto 18) &
  n17(17 downto 17);
process (clock_c) begin
  if rising_edge(clock_c) then
    if i5 = "1" then
      n19 <= "000000000000000000";
    elsif i4 = "1" then
      n19 <= n18;
    end if;
  end if;
end process;
n20 <= n16 - n19;
process (clock_c) begin
  if rising_edge(clock_c) then
    if i5 = "1" then
      n21 <= "000000000000000000";
    elsif i4 = "1" then
      n21 <= n20;
    end if;
  end if;
end process;
n22 <= unsigned(signed(n5) * signed(n13));
n23 <= n22(34 downto 34) &
  n22(33 downto 33) &
  n22(32 downto 32) &
  n22(31 downto 31) &
  n22(30 downto 30) &
  n22(29 downto 29) &
  n22(28 downto 28) &
  n22(27 downto 27) &
  n22(26 downto 26) &
  n22(25 downto 25) &
  n22(24 downto 24) &
  n22(23 downto 23) &
  n22(22 downto 22) &
  n22(21 downto 21) &
  n22(20 downto 20) &
  n22(19 downto 19) &
  n22(18 downto 18) &
  n22(17 downto 17);
process (clock_c) begin
  if rising_edge(clock_c) then
    if i5 = "1" then
      n24 <= "000000000000000000";
    elsif i4 = "1" then
      n24 <= n23;
    end if;
  end if;
end process;
n25 <= unsigned(signed(n6) * signed(n12));
n26 <= n25(34 downto 34) &
  n25(33 downto 33) &
  n25(32 downto 32) &
  n25(31 downto 31) &
  n25(30 downto 30) &
  n25(29 downto 29) &
  n25(28 downto 28) &
  n25(27 downto 27) &
  n25(26 downto 26) &
  n25(25 downto 25) &
  n25(24 downto 24) &
  n25(23 downto 23) &
  n25(22 downto 22) &
  n25(21 downto 21) &
  n25(20 downto 20) &
  n25(19 downto 19) &
  n25(18 downto 18) &
  n25(17 downto 17);
process (clock_c) begin
  if rising_edge(clock_c) then
    if i5 = "1" then
      n27 <= "000000000000000000";
    elsif i4 = "1" then
      n27 <= n26;
    end if;
  end if;
end process;
n28 <= n24 + n27;
process (clock_c) begin
  if rising_edge(clock_c) then
    if i5 = "1" then
      n29 <= "000000000000000000";
    elsif i4 = "1" then
      n29 <= n28;
    end if;
  end if;
end process;
n30 <= n8 + n21;
n31 <= n10 + n29;
n32 <= n30 & n31;
process (clock_c) begin
  if rising_edge(clock_c) then
    if i5 = "1" then
      n33 <= "000000000000000000000000000000000000";
    elsif i4 = "1" then
      n33 <= n32;
    end if;
  end if;
end process;
n34 <= n8 - n21;
n35 <= n10 - n29;
n36 <= n34 & n35;
process (clock_c) begin
  if rising_edge(clock_c) then
    if i5 = "1" then
      n37 <= "000000000000000000000000000000000000";
    elsif i4 = "1" then
      n37 <= n36;
    end if;
  end if;
end process;
o2 <= n37;
o1 <= n33;
end architecture rtl;

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
entity cf_fft_4096_18_23 is
port (
clock_c : in std_logic;
i1 : in  unsigned(0 downto 0);
i2 : in  unsigned(35 downto 0);
i3 : in  unsigned(35 downto 0);
i4 : in  unsigned(0 downto 0);
i5 : in  unsigned(0 downto 0);
o1 : out unsigned(0 downto 0);
o2 : out unsigned(35 downto 0);
o3 : out unsigned(35 downto 0));
end entity cf_fft_4096_18_23;
architecture rtl of cf_fft_4096_18_23 is
signal n1 : unsigned(9 downto 0);
signal n2 : unsigned(71 downto 0);
signal n3 : unsigned(0 downto 0) := "0";
signal n4 : unsigned(0 downto 0) := "0";
signal n5 : unsigned(0 downto 0) := "0";
signal n6 : unsigned(0 downto 0) := "0";
signal n7 : unsigned(9 downto 0);
signal n8 : unsigned(9 downto 0) := "0000000000";
signal n9 : unsigned(9 downto 0) := "0000000000";
signal n10 : unsigned(9 downto 0) := "0000000000";
signal n11 : unsigned(9 downto 0) := "0000000000";
signal n12 : unsigned(0 downto 0);
signal n13 : unsigned(0 downto 0) := "0";
signal n14 : unsigned(0 downto 0) := "0";
signal n15 : unsigned(0 downto 0) := "0";
signal n16 : unsigned(0 downto 0) := "0";
signal n17 : unsigned(0 downto 0);
signal n18 : unsigned(1 downto 0);
signal n19 : unsigned(35 downto 0);
signal n20 : unsigned(35 downto 0);
signal n21 : unsigned(35 downto 0);
signal n22 : unsigned(35 downto 0);
signal n23 : unsigned(35 downto 0);
signal n24 : unsigned(35 downto 0);
signal s25_1 : unsigned(35 downto 0);
signal s25_2 : unsigned(35 downto 0);
signal s26_1 : unsigned(0 downto 0);
signal s27_1 : unsigned(71 downto 0);
signal s28_1 : unsigned(0 downto 0);
signal s28_2 : unsigned(0 downto 0);
signal s28_3 : unsigned(71 downto 0);
signal s29_1 : unsigned(10 downto 0);
signal s29_2 : unsigned(0 downto 0);
component cf_fft_4096_18_24 is
port (
clock_c : in std_logic;
i1 : in  unsigned(35 downto 0);
i2 : in  unsigned(35 downto 0);
i3 : in  unsigned(9 downto 0);
i4 : in  unsigned(0 downto 0);
i5 : in  unsigned(0 downto 0);
o1 : out unsigned(35 downto 0);
o2 : out unsigned(35 downto 0));
end component cf_fft_4096_18_24;
component cf_fft_4096_18_37 is
port (
clock_c : in std_logic;
i1 : in  unsigned(1 downto 0);
i2 : in  unsigned(0 downto 0);
i3 : in  unsigned(0 downto 0);
o1 : out unsigned(0 downto 0));
end component cf_fft_4096_18_37;
component cf_fft_4096_18_33 is
port (
clock_c : in std_logic;
i1 : in  unsigned(71 downto 0);
i2 : in  unsigned(0 downto 0);
i3 : in  unsigned(9 downto 0);
i4 : in  unsigned(0 downto 0);
i5 : in  unsigned(0 downto 0);
i6 : in  unsigned(0 downto 0);
o1 : out unsigned(71 downto 0));
end component cf_fft_4096_18_33;
component cf_fft_4096_18_32 is
port (
clock_c : in std_logic;
i1 : in  unsigned(71 downto 0);
i2 : in  unsigned(0 downto 0);
i3 : in  unsigned(9 downto 0);
i4 : in  unsigned(0 downto 0);
i5 : in  unsigned(0 downto 0);
i6 : in  unsigned(0 downto 0);
o1 : out unsigned(0 downto 0);
o2 : out unsigned(0 downto 0);
o3 : out unsigned(71 downto 0));
end component cf_fft_4096_18_32;
component cf_fft_4096_18_28 is
port (
clock_c : in std_logic;
i1 : in  unsigned(0 downto 0);
i2 : in  unsigned(0 downto 0);
i3 : in  unsigned(0 downto 0);
o1 : out unsigned(10 downto 0);
o2 : out unsigned(0 downto 0));
end component cf_fft_4096_18_28;
begin
n1 <= s29_1(10 downto 10) &
  s29_1(9 downto 9) &
  s29_1(8 downto 8) &
  s29_1(7 downto 7) &
  s29_1(6 downto 6) &
  s29_1(5 downto 5) &
  s29_1(4 downto 4) &
  s29_1(3 downto 3) &
  s29_1(2 downto 2) &
  s29_1(1 downto 1);
n2 <= s25_1 & s25_2;
process (clock_c) begin
  if rising_edge(clock_c) then
    if i5 = "1" then
      n3 <= "0";
    elsif i4 = "1" then
      n3 <= s29_2;
    end if;
  end if;
end process;
process (clock_c) begin
  if rising_edge(clock_c) then
    if i5 = "1" then
      n4 <= "0";
    elsif i4 = "1" then
      n4 <= n3;
    end if;
  end if;
end process;
process (clock_c) begin
  if rising_edge(clock_c) then
    if i5 = "1" then
      n5 <= "0";
    elsif i4 = "1" then
      n5 <= n4;
    end if;
  end if;
end process;
process (clock_c) begin
  if rising_edge(clock_c) then
    if i5 = "1" then
      n6 <= "0";
    elsif i4 = "1" then
      n6 <= n5;
    end if;
  end if;
end process;
n7 <= s29_1(10 downto 10) &
  s29_1(9 downto 9) &
  s29_1(8 downto 8) &
  s29_1(7 downto 7) &
  s29_1(6 downto 6) &
  s29_1(5 downto 5) &
  s29_1(4 downto 4) &
  s29_1(3 downto 3) &
  s29_1(2 downto 2) &
  s29_1(1 downto 1);
process (clock_c) begin
  if rising_edge(clock_c) then
    if i5 = "1" then
      n8 <= "0000000000";
    elsif i4 = "1" then
      n8 <= n7;
    end if;
  end if;
end process;
process (clock_c) begin
  if rising_edge(clock_c) then
    if i5 = "1" then
      n9 <= "0000000000";
    elsif i4 = "1" then
      n9 <= n8;
    end if;
  end if;
end process;
process (clock_c) begin
  if rising_edge(clock_c) then
    if i5 = "1" then
      n10 <= "0000000000";
    elsif i4 = "1" then
      n10 <= n9;
    end if;
  end if;
end process;
process (clock_c) begin
  if rising_edge(clock_c) then
    if i5 = "1" then
      n11 <= "0000000000";
    elsif i4 = "1" then
      n11 <= n10;
    end if;
  end if;
end process;
n12 <= s29_1(0 downto 0);
process (clock_c) begin
  if rising_edge(clock_c) then
    if i5 = "1" then
      n13 <= "0";
    elsif i4 = "1" then
      n13 <= n12;
    end if;
  end if;
end process;
process (clock_c) begin
  if rising_edge(clock_c) then
    if i5 = "1" then
      n14 <= "0";
    elsif i4 = "1" then
      n14 <= n13;
    end if;
  end if;
end process;
process (clock_c) begin
  if rising_edge(clock_c) then
    if i5 = "1" then
      n15 <= "0";
    elsif i4 = "1" then
      n15 <= n14;
    end if;
  end if;
end process;
process (clock_c) begin
  if rising_edge(clock_c) then
    if i5 = "1" then
      n16 <= "0";
    elsif i4 = "1" then
      n16 <= n15;
    end if;
  end if;
end process;
n17 <= not n16;
n18 <= s28_2 & s28_1;
n19 <= s28_3(71 downto 71) &
  s28_3(70 downto 70) &
  s28_3(69 downto 69) &
  s28_3(68 downto 68) &
  s28_3(67 downto 67) &
  s28_3(66 downto 66) &
  s28_3(65 downto 65) &
  s28_3(64 downto 64) &
  s28_3(63 downto 63) &
  s28_3(62 downto 62) &
  s28_3(61 downto 61) &
  s28_3(60 downto 60) &
  s28_3(59 downto 59) &
  s28_3(58 downto 58) &
  s28_3(57 downto 57) &
  s28_3(56 downto 56) &
  s28_3(55 downto 55) &
  s28_3(54 downto 54) &
  s28_3(53 downto 53) &
  s28_3(52 downto 52) &
  s28_3(51 downto 51) &
  s28_3(50 downto 50) &
  s28_3(49 downto 49) &
  s28_3(48 downto 48) &
  s28_3(47 downto 47) &
  s28_3(46 downto 46) &
  s28_3(45 downto 45) &
  s28_3(44 downto 44) &
  s28_3(43 downto 43) &
  s28_3(42 downto 42) &
  s28_3(41 downto 41) &
  s28_3(40 downto 40) &
  s28_3(39 downto 39) &
  s28_3(38 downto 38) &
  s28_3(37 downto 37) &
  s28_3(36 downto 36);
n20 <= s28_3(35 downto 35) &
  s28_3(34 downto 34) &
  s28_3(33 downto 33) &
  s28_3(32 downto 32) &
  s28_3(31 downto 31) &
  s28_3(30 downto 30) &
  s28_3(29 downto 29) &
  s28_3(28 downto 28) &
  s28_3(27 downto 27) &
  s28_3(26 downto 26) &
  s28_3(25 downto 25) &
  s28_3(24 downto 24) &
  s28_3(23 downto 23) &
  s28_3(22 downto 22) &
  s28_3(21 downto 21) &
  s28_3(20 downto 20) &
  s28_3(19 downto 19) &
  s28_3(18 downto 18) &
  s28_3(17 downto 17) &
  s28_3(16 downto 16) &
  s28_3(15 downto 15) &
  s28_3(14 downto 14) &
  s28_3(13 downto 13) &
  s28_3(12 downto 12) &
  s28_3(11 downto 11) &
  s28_3(10 downto 10) &
  s28_3(9 downto 9) &
  s28_3(8 downto 8) &
  s28_3(7 downto 7) &
  s28_3(6 downto 6) &
  s28_3(5 downto 5) &
  s28_3(4 downto 4) &
  s28_3(3 downto 3) &
  s28_3(2 downto 2) &
  s28_3(1 downto 1) &
  s28_3(0 downto 0);
n21 <= s27_1(71 downto 71) &
  s27_1(70 downto 70) &
  s27_1(69 downto 69) &
  s27_1(68 downto 68) &
  s27_1(67 downto 67) &
  s27_1(66 downto 66) &
  s27_1(65 downto 65) &
  s27_1(64 downto 64) &
  s27_1(63 downto 63) &
  s27_1(62 downto 62) &
  s27_1(61 downto 61) &
  s27_1(60 downto 60) &
  s27_1(59 downto 59) &
  s27_1(58 downto 58) &
  s27_1(57 downto 57) &
  s27_1(56 downto 56) &
  s27_1(55 downto 55) &
  s27_1(54 downto 54) &
  s27_1(53 downto 53) &
  s27_1(52 downto 52) &
  s27_1(51 downto 51) &
  s27_1(50 downto 50) &
  s27_1(49 downto 49) &
  s27_1(48 downto 48) &
  s27_1(47 downto 47) &
  s27_1(46 downto 46) &
  s27_1(45 downto 45) &
  s27_1(44 downto 44) &
  s27_1(43 downto 43) &
  s27_1(42 downto 42) &
  s27_1(41 downto 41) &
  s27_1(40 downto 40) &
  s27_1(39 downto 39) &
  s27_1(38 downto 38) &
  s27_1(37 downto 37) &
  s27_1(36 downto 36);
n22 <= s27_1(35 downto 35) &
  s27_1(34 downto 34) &
  s27_1(33 downto 33) &
  s27_1(32 downto 32) &
  s27_1(31 downto 31) &
  s27_1(30 downto 30) &
  s27_1(29 downto 29) &
  s27_1(28 downto 28) &
  s27_1(27 downto 27) &
  s27_1(26 downto 26) &
  s27_1(25 downto 25) &
  s27_1(24 downto 24) &
  s27_1(23 downto 23) &
  s27_1(22 downto 22) &
  s27_1(21 downto 21) &
  s27_1(20 downto 20) &
  s27_1(19 downto 19) &
  s27_1(18 downto 18) &
  s27_1(17 downto 17) &
  s27_1(16 downto 16) &
  s27_1(15 downto 15) &
  s27_1(14 downto 14) &
  s27_1(13 downto 13) &
  s27_1(12 downto 12) &
  s27_1(11 downto 11) &
  s27_1(10 downto 10) &
  s27_1(9 downto 9) &
  s27_1(8 downto 8) &
  s27_1(7 downto 7) &
  s27_1(6 downto 6) &
  s27_1(5 downto 5) &
  s27_1(4 downto 4) &
  s27_1(3 downto 3) &
  s27_1(2 downto 2) &
  s27_1(1 downto 1) &
  s27_1(0 downto 0);
n23 <= n20 when s26_1 = "1" else n19;
n24 <= n22 when s26_1 = "1" else n21;
s25 : cf_fft_4096_18_24 port map (clock_c, i2, i3, n1, i4, i5, s25_1, s25_2);
s26 : cf_fft_4096_18_37 port map (clock_c, n18, i4, i5, s26_1);
s27 : cf_fft_4096_18_33 port map (clock_c, n2, n6, n11, n16, i4, i5, s27_1);
s28 : cf_fft_4096_18_32 port map (clock_c, n2, n6, n11, n17, i4, i5, s28_1, s28_2, s28_3);
s29 : cf_fft_4096_18_28 port map (clock_c, i1, i4, i5, s29_1, s29_2);
o3 <= n24;
o2 <= n23;
o1 <= s28_1;
end architecture rtl;

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
entity cf_fft_4096_18_22 is
port (
clock_c : in std_logic;
i1 : in  unsigned(35 downto 0);
i2 : in  unsigned(35 downto 0);
i3 : in  unsigned(8 downto 0);
i4 : in  unsigned(0 downto 0);
i5 : in  unsigned(0 downto 0);
o1 : out unsigned(35 downto 0);
o2 : out unsigned(35 downto 0));
end entity cf_fft_4096_18_22;
architecture rtl of cf_fft_4096_18_22 is
signal n1 : unsigned(35 downto 0) := "000000000000000000000000000000000000";
signal n2 : unsigned(17 downto 0);
signal n3 : unsigned(17 downto 0);
signal n4 : unsigned(35 downto 0) := "000000000000000000000000000000000000";
signal n5 : unsigned(17 downto 0);
signal n6 : unsigned(17 downto 0);
signal n7 : unsigned(17 downto 0) := "000000000000000000";
signal n8 : unsigned(17 downto 0) := "000000000000000000";
signal n9 : unsigned(17 downto 0) := "000000000000000000";
signal n10 : unsigned(17 downto 0) := "000000000000000000";
signal n11 : unsigned(35 downto 0) := "000000000000000000000000000000000000";
signal n12 : unsigned(17 downto 0);
signal n13 : unsigned(17 downto 0);
signal n14 : unsigned(35 downto 0);
signal n15 : unsigned(17 downto 0);
signal n16 : unsigned(17 downto 0) := "000000000000000000";
signal n17 : unsigned(35 downto 0);
signal n18 : unsigned(17 downto 0);
signal n19 : unsigned(17 downto 0) := "000000000000000000";
signal n20 : unsigned(17 downto 0);
signal n21 : unsigned(17 downto 0) := "000000000000000000";
signal n22 : unsigned(35 downto 0);
signal n23 : unsigned(17 downto 0);
signal n24 : unsigned(17 downto 0) := "000000000000000000";
signal n25 : unsigned(35 downto 0);
signal n26 : unsigned(17 downto 0);
signal n27 : unsigned(17 downto 0) := "000000000000000000";
signal n28 : unsigned(17 downto 0);
signal n29 : unsigned(17 downto 0) := "000000000000000000";
signal n30 : unsigned(17 downto 0);
signal n31 : unsigned(17 downto 0);
signal n32 : unsigned(35 downto 0);
signal n33 : unsigned(35 downto 0) := "000000000000000000000000000000000000";
signal n34 : unsigned(17 downto 0);
signal n35 : unsigned(17 downto 0);
signal n36 : unsigned(35 downto 0);
signal n37 : unsigned(35 downto 0) := "000000000000000000000000000000000000";
begin
process (clock_c) begin
  if rising_edge(clock_c) then
    if i5 = "1" then
      n1 <= "000000000000000000000000000000000000";
    elsif i4 = "1" then
      n1 <= i1;
    end if;
  end if;
end process;
n2 <= n1(35 downto 35) &
  n1(34 downto 34) &
  n1(33 downto 33) &
  n1(32 downto 32) &
  n1(31 downto 31) &
  n1(30 downto 30) &
  n1(29 downto 29) &
  n1(28 downto 28) &
  n1(27 downto 27) &
  n1(26 downto 26) &
  n1(25 downto 25) &
  n1(24 downto 24) &
  n1(23 downto 23) &
  n1(22 downto 22) &
  n1(21 downto 21) &
  n1(20 downto 20) &
  n1(19 downto 19) &
  n1(18 downto 18);
n3 <= n1(17 downto 17) &
  n1(16 downto 16) &
  n1(15 downto 15) &
  n1(14 downto 14) &
  n1(13 downto 13) &
  n1(12 downto 12) &
  n1(11 downto 11) &
  n1(10 downto 10) &
  n1(9 downto 9) &
  n1(8 downto 8) &
  n1(7 downto 7) &
  n1(6 downto 6) &
  n1(5 downto 5) &
  n1(4 downto 4) &
  n1(3 downto 3) &
  n1(2 downto 2) &
  n1(1 downto 1) &
  n1(0 downto 0);
process (clock_c) begin
  if rising_edge(clock_c) then
    if i5 = "1" then
      n4 <= "000000000000000000000000000000000000";
    elsif i4 = "1" then
      n4 <= i2;
    end if;
  end if;
end process;
n5 <= n4(35 downto 35) &
  n4(34 downto 34) &
  n4(33 downto 33) &
  n4(32 downto 32) &
  n4(31 downto 31) &
  n4(30 downto 30) &
  n4(29 downto 29) &
  n4(28 downto 28) &
  n4(27 downto 27) &
  n4(26 downto 26) &
  n4(25 downto 25) &
  n4(24 downto 24) &
  n4(23 downto 23) &
  n4(22 downto 22) &
  n4(21 downto 21) &
  n4(20 downto 20) &
  n4(19 downto 19) &
  n4(18 downto 18);
n6 <= n4(17 downto 17) &
  n4(16 downto 16) &
  n4(15 downto 15) &
  n4(14 downto 14) &
  n4(13 downto 13) &
  n4(12 downto 12) &
  n4(11 downto 11) &
  n4(10 downto 10) &
  n4(9 downto 9) &
  n4(8 downto 8) &
  n4(7 downto 7) &
  n4(6 downto 6) &
  n4(5 downto 5) &
  n4(4 downto 4) &
  n4(3 downto 3) &
  n4(2 downto 2) &
  n4(1 downto 1) &
  n4(0 downto 0);
process (clock_c) begin
  if rising_edge(clock_c) then
    if i5 = "1" then
      n7 <= "000000000000000000";
    elsif i4 = "1" then
      n7 <= n2;
    end if;
  end if;
end process;
process (clock_c) begin
  if rising_edge(clock_c) then
    if i5 = "1" then
      n8 <= "000000000000000000";
    elsif i4 = "1" then
      n8 <= n7;
    end if;
  end if;
end process;
process (clock_c) begin
  if rising_edge(clock_c) then
    if i5 = "1" then
      n9 <= "000000000000000000";
    elsif i4 = "1" then
      n9 <= n3;
    end if;
  end if;
end process;
process (clock_c) begin
  if rising_edge(clock_c) then
    if i5 = "1" then
      n10 <= "000000000000000000";
    elsif i4 = "1" then
      n10 <= n9;
    end if;
  end if;
end process;
process (clock_c) begin
  if rising_edge(clock_c) then 
    if i4 = "1" then
      case i3 is
        when "000000000" => n11 <= "011111111111111111000000000000000000";
        when "000000001" => n11 <= "011111111111111101111111110011011011";
        when "000000010" => n11 <= "011111111111110110111111100110110111";
        when "000000011" => n11 <= "011111111111101001111111011010010011";
        when "000000100" => n11 <= "011111111111011000111111001101101111";
        when "000000101" => n11 <= "011111111111000010111111000001001011";
        when "000000110" => n11 <= "011111111110100111111110110100100111";
        when "000000111" => n11 <= "011111111110000111111110101000000011";
        when "000001000" => n11 <= "011111111101100010111110011011100000";
        when "000001001" => n11 <= "011111111100111000111110001110111101";
        when "000001010" => n11 <= "011111111100001001111110000010011010";
        when "000001011" => n11 <= "011111111011010101111101110101110111";
        when "000001100" => n11 <= "011111111010011100111101101001010101";
        when "000001101" => n11 <= "011111111001011111111101011100110011";
        when "000001110" => n11 <= "011111111000011100111101010000010010";
        when "000001111" => n11 <= "011111110111010101111101000011110001";
        when "000010000" => n11 <= "011111110110001000111100110111010000";
        when "000010001" => n11 <= "011111110100110111111100101010110000";
        when "000010010" => n11 <= "011111110011100001111100011110010000";
        when "000010011" => n11 <= "011111110010000110111100010001110001";
        when "000010100" => n11 <= "011111110000100110111100000101010011";
        when "000010101" => n11 <= "011111101111000001111011111000110101";
        when "000010110" => n11 <= "011111101101010111111011101100011000";
        when "000010111" => n11 <= "011111101011101000111011011111111011";
        when "000011000" => n11 <= "011111101001110101111011010011011111";
        when "000011001" => n11 <= "011111100111111100111011000111000100";
        when "000011010" => n11 <= "011111100101111111111010111010101010";
        when "000011011" => n11 <= "011111100011111101111010101110010000";
        when "000011100" => n11 <= "011111100001110110111010100001110111";
        when "000011101" => n11 <= "011111011111101010111010010101011111";
        when "000011110" => n11 <= "011111011101011001111010001001001000";
        when "000011111" => n11 <= "011111011011000011111001111100110010";
        when "000100000" => n11 <= "011111011000101001111001110000011101";
        when "000100001" => n11 <= "011111010110001010111001100100001000";
        when "000100010" => n11 <= "011111010011100110111001010111110101";
        when "000100011" => n11 <= "011111010000111101111001001011100011";
        when "000100100" => n11 <= "011111001110001111111000111111010001";
        when "000100101" => n11 <= "011111001011011100111000110011000001";
        when "000100110" => n11 <= "011111001000100101111000100110110010";
        when "000100111" => n11 <= "011111000101101000111000011010100100";
        when "000101000" => n11 <= "011111000010100111111000001110011000";
        when "000101001" => n11 <= "011110111111100010111000000010001100";
        when "000101010" => n11 <= "011110111100010111110111110110000010";
        when "000101011" => n11 <= "011110111001001000110111101001111001";
        when "000101100" => n11 <= "011110110101110100110111011101110001";
        when "000101101" => n11 <= "011110110010011011110111010001101010";
        when "000101110" => n11 <= "011110101110111101110111000101100101";
        when "000101111" => n11 <= "011110101011011011110110111001100010";
        when "000110000" => n11 <= "011110100111110100110110101101011111";
        when "000110001" => n11 <= "011110100100001000110110100001011110";
        when "000110010" => n11 <= "011110100000010111110110010101011111";
        when "000110011" => n11 <= "011110011100100010110110001001100001";
        when "000110100" => n11 <= "011110011000101000110101111101100101";
        when "000110101" => n11 <= "011110010100101001110101110001101010";
        when "000110110" => n11 <= "011110010000100110110101100101110000";
        when "000110111" => n11 <= "011110001100011110110101011001111001";
        when "000111000" => n11 <= "011110001000010010110101001110000011";
        when "000111001" => n11 <= "011110000100000000110101000010001110";
        when "000111010" => n11 <= "011101111111101010110100110110011100";
        when "000111011" => n11 <= "011101111011010000110100101010101011";
        when "000111100" => n11 <= "011101110110110001110100011110111011";
        when "000111101" => n11 <= "011101110010001101110100010011001110";
        when "000111110" => n11 <= "011101101101100101110100000111100010";
        when "000111111" => n11 <= "011101101000111000110011111011111000";
        when "001000000" => n11 <= "011101100100000110110011110000010000";
        when "001000001" => n11 <= "011101011111010000110011100100101010";
        when "001000010" => n11 <= "011101011010010110110011011001000110";
        when "001000011" => n11 <= "011101010101010110110011001101100100";
        when "001000100" => n11 <= "011101010000010011110011000010000100";
        when "001000101" => n11 <= "011101001011001011110010110110100101";
        when "001000110" => n11 <= "011101000101111110110010101011001001";
        when "001000111" => n11 <= "011101000000101101110010011111101111";
        when "001001000" => n11 <= "011100111011010111110010010100010111";
        when "001001001" => n11 <= "011100110101111101110010001001000001";
        when "001001010" => n11 <= "011100110000011111110001111101101101";
        when "001001011" => n11 <= "011100101010111100110001110010011100";
        when "001001100" => n11 <= "011100100101010100110001100111001100";
        when "001001101" => n11 <= "011100011111101000110001011011111111";
        when "001001110" => n11 <= "011100011001111000110001010000110100";
        when "001001111" => n11 <= "011100010100000100110001000101101011";
        when "001010000" => n11 <= "011100001110001011110000111010100101";
        when "001010001" => n11 <= "011100001000001101110000101111100000";
        when "001010010" => n11 <= "011100000010001100110000100100011111";
        when "001010011" => n11 <= "011011111100000110110000011001011111";
        when "001010100" => n11 <= "011011110101111100110000001110100010";
        when "001010101" => n11 <= "011011101111101101110000000011101000";
        when "001010110" => n11 <= "011011101001011010101111111000110000";
        when "001010111" => n11 <= "011011100011000011101111101101111010";
        when "001011000" => n11 <= "011011011100101000101111100011000111";
        when "001011001" => n11 <= "011011010110001000101111011000010110";
        when "001011010" => n11 <= "011011001111100100101111001101101000";
        when "001011011" => n11 <= "011011001000111100101111000010111101";
        when "001011100" => n11 <= "011011000010010000101110111000010100";
        when "001011101" => n11 <= "011010111011100000101110101101101110";
        when "001011110" => n11 <= "011010110100101011101110100011001011";
        when "001011111" => n11 <= "011010101101110011101110011000101010";
        when "001100000" => n11 <= "011010100110110110101110001110001100";
        when "001100001" => n11 <= "011010011111110101101110000011110000";
        when "001100010" => n11 <= "011010011000110000101101111001011000";
        when "001100011" => n11 <= "011010010001100111101101101111000010";
        when "001100100" => n11 <= "011010001010011010101101100100101111";
        when "001100101" => n11 <= "011010000011001001101101011010011111";
        when "001100110" => n11 <= "011001111011110100101101010000010010";
        when "001100111" => n11 <= "011001110100011011101101000110000111";
        when "001101000" => n11 <= "011001101100111110101100111100000000";
        when "001101001" => n11 <= "011001100101011100101100110001111011";
        when "001101010" => n11 <= "011001011101110111101100100111111010";
        when "001101011" => n11 <= "011001010110001110101100011101111011";
        when "001101100" => n11 <= "011001001110100010101100010100000000";
        when "001101101" => n11 <= "011001000110110001101100001010000111";
        when "001101110" => n11 <= "011000111110111100101100000000010010";
        when "001101111" => n11 <= "011000110111000100101011110110100000";
        when "001110000" => n11 <= "011000101111001000101011101100110000";
        when "001110001" => n11 <= "011000100111000111101011100011000100";
        when "001110010" => n11 <= "011000011111000100101011011001011011";
        when "001110011" => n11 <= "011000010110111100101011001111110101";
        when "001110100" => n11 <= "011000001110110000101011000110010011";
        when "001110101" => n11 <= "011000000110100001101010111100110011";
        when "001110110" => n11 <= "010111111110001110101010110011010111";
        when "001110111" => n11 <= "010111110101111000101010101001111110";
        when "001111000" => n11 <= "010111101101011101101010100000101001";
        when "001111001" => n11 <= "010111100101000000101010010111010111";
        when "001111010" => n11 <= "010111011100011110101010001110001000";
        when "001111011" => n11 <= "010111010011111001101010000100111100";
        when "001111100" => n11 <= "010111001011010000101001111011110100";
        when "001111101" => n11 <= "010111000010100100101001110010101111";
        when "001111110" => n11 <= "010110111001110100101001101001101110";
        when "001111111" => n11 <= "010110110001000000101001100000110000";
        when "010000000" => n11 <= "010110101000001001101001010111110110";
        when "010000001" => n11 <= "010110011111001111101001001110111111";
        when "010000010" => n11 <= "010110010110010001101001000110001011";
        when "010000011" => n11 <= "010110001101010000101000111101011011";
        when "010000100" => n11 <= "010110000100001011101000110100101111";
        when "010000101" => n11 <= "010101111011000011101000101100000110";
        when "010000110" => n11 <= "010101110001110111101000100011100001";
        when "010000111" => n11 <= "010101101000101000101000011010111111";
        when "010001000" => n11 <= "010101011111010110101000010010100010";
        when "010001001" => n11 <= "010101010110000001101000001010000111";
        when "010001010" => n11 <= "010101001100101000101000000001110001";
        when "010001011" => n11 <= "010101000011001100100111111001011110";
        when "010001100" => n11 <= "010100111001101100100111110001001111";
        when "010001101" => n11 <= "010100110000001010100111101001000011";
        when "010001110" => n11 <= "010100100110100100100111100000111011";
        when "010001111" => n11 <= "010100011100111011100111011000111000";
        when "010010000" => n11 <= "010100010011001111100111010000110111";
        when "010010001" => n11 <= "010100001001011111100111001000111011";
        when "010010010" => n11 <= "010011111111101101100111000001000011";
        when "010010011" => n11 <= "010011110101111000100110111001001110";
        when "010010100" => n11 <= "010011101011111111100110110001011101";
        when "010010101" => n11 <= "010011100010000100100110101001110001";
        when "010010110" => n11 <= "010011011000000101100110100010001000";
        when "010010111" => n11 <= "010011001110000100100110011010100011";
        when "010011000" => n11 <= "010011000011111111100110010011000001";
        when "010011001" => n11 <= "010010111001111000100110001011100100";
        when "010011010" => n11 <= "010010101111101101100110000100001011";
        when "010011011" => n11 <= "010010100101100000100101111100110110";
        when "010011100" => n11 <= "010010011011010000100101110101100101";
        when "010011101" => n11 <= "010010010000111101100101101110011000";
        when "010011110" => n11 <= "010010000110100111100101100111001111";
        when "010011111" => n11 <= "010001111100001111100101100000001010";
        when "010100000" => n11 <= "010001110001110011100101011001001001";
        when "010100001" => n11 <= "010001100111010101100101010010001100";
        when "010100010" => n11 <= "010001011100110100100101001011010100";
        when "010100011" => n11 <= "010001010010010001100101000100011111";
        when "010100100" => n11 <= "010001000111101011100100111101101111";
        when "010100101" => n11 <= "010000111101000010100100110111000011";
        when "010100110" => n11 <= "010000110010010111100100110000011011";
        when "010100111" => n11 <= "010000100111101001100100101001110111";
        when "010101000" => n11 <= "010000011100111000100100100011010111";
        when "010101001" => n11 <= "010000010010000101100100011100111100";
        when "010101010" => n11 <= "010000000111001111100100010110100101";
        when "010101011" => n11 <= "001111111100010111100100010000010010";
        when "010101100" => n11 <= "001111110001011101100100001010000011";
        when "010101101" => n11 <= "001111100110100000100100000011111001";
        when "010101110" => n11 <= "001111011011100000100011111101110011";
        when "010101111" => n11 <= "001111010000011111100011110111110010";
        when "010110000" => n11 <= "001111000101011010100011110001110100";
        when "010110001" => n11 <= "001110111010010100100011101011111011";
        when "010110010" => n11 <= "001110101111001011100011100110000111";
        when "010110011" => n11 <= "001110100100000000100011100000010111";
        when "010110100" => n11 <= "001110011000110011100011011010101011";
        when "010110101" => n11 <= "001110001101100011100011010101000011";
        when "010110110" => n11 <= "001110000010010010100011001111100000";
        when "010110111" => n11 <= "001101110110111110100011001010000010";
        when "010111000" => n11 <= "001101101011101000100011000100101000";
        when "010111001" => n11 <= "001101100000010000100010111111010010";
        when "010111010" => n11 <= "001101010100110110100010111010000001";
        when "010111011" => n11 <= "001101001001011010100010110100110100";
        when "010111100" => n11 <= "001100111101111011100010101111101100";
        when "010111101" => n11 <= "001100110010011011100010101010101001";
        when "010111110" => n11 <= "001100100110111001100010100101101001";
        when "010111111" => n11 <= "001100011011010101100010100000101111";
        when "011000000" => n11 <= "001100001111101111100010011011111001";
        when "011000001" => n11 <= "001100000100000111100010010111000111";
        when "011000010" => n11 <= "001011111000011101100010010010011010";
        when "011000011" => n11 <= "001011101100110001100010001101110010";
        when "011000100" => n11 <= "001011100001000100100010001001001110";
        when "011000101" => n11 <= "001011010101010100100010000100101111";
        when "011000110" => n11 <= "001011001001100011100010000000010101";
        when "011000111" => n11 <= "001010111101110001100001111011111111";
        when "011001000" => n11 <= "001010110001111100100001110111101101";
        when "011001001" => n11 <= "001010100110000110100001110011100001";
        when "011001010" => n11 <= "001010011010001111100001101111011001";
        when "011001011" => n11 <= "001010001110010101100001101011010110";
        when "011001100" => n11 <= "001010000010011010100001100111010111";
        when "011001101" => n11 <= "001001110110011110100001100011011101";
        when "011001110" => n11 <= "001001101010100000100001011111101000";
        when "011001111" => n11 <= "001001011110100001100001011011110111";
        when "011010000" => n11 <= "001001010010100000100001011000001011";
        when "011010001" => n11 <= "001001000110011101100001010100100100";
        when "011010010" => n11 <= "001000111010011010100001010001000010";
        when "011010011" => n11 <= "001000101110010101100001001101100100";
        when "011010100" => n11 <= "001000100010001110100001001010001011";
        when "011010101" => n11 <= "001000010110000110100001000110110111";
        when "011010110" => n11 <= "001000001001111101100001000011101000";
        when "011010111" => n11 <= "000111111101110011100001000000011101";
        when "011011000" => n11 <= "000111110001100111100000111101011000";
        when "011011001" => n11 <= "000111100101011011100000111010010111";
        when "011011010" => n11 <= "000111011001001101100000110111011010";
        when "011011011" => n11 <= "000111001100111110100000110100100011";
        when "011011100" => n11 <= "000111000000101110100000110001110000";
        when "011011101" => n11 <= "000110110100011100100000101111000010";
        when "011011110" => n11 <= "000110101000001010100000101100011001";
        when "011011111" => n11 <= "000110011011110111100000101001110101";
        when "011100000" => n11 <= "000110001111100010100000100111010110";
        when "011100001" => n11 <= "000110000011001101100000100100111100";
        when "011100010" => n11 <= "000101110110110111100000100010100110";
        when "011100011" => n11 <= "000101101010100000100000100000010101";
        when "011100100" => n11 <= "000101011110001000100000011110001001";
        when "011100101" => n11 <= "000101010001101111100000011100000010";
        when "011100110" => n11 <= "000101000101010101100000011010000000";
        when "011100111" => n11 <= "000100111000111011100000011000000011";
        when "011101000" => n11 <= "000100101100100000100000010110001010";
        when "011101001" => n11 <= "000100100000000100100000010100010111";
        when "011101010" => n11 <= "000100010011100111100000010010101000";
        when "011101011" => n11 <= "000100000111001010100000010000111110";
        when "011101100" => n11 <= "000011111010101100100000001111011001";
        when "011101101" => n11 <= "000011101110001110100000001101111001";
        when "011101110" => n11 <= "000011100001101111100000001100011110";
        when "011101111" => n11 <= "000011010101001111100000001011001000";
        when "011110000" => n11 <= "000011001000101111100000001001110111";
        when "011110001" => n11 <= "000010111100001110100000001000101010";
        when "011110010" => n11 <= "000010101111101101100000000111100011";
        when "011110011" => n11 <= "000010100011001100100000000110100000";
        when "011110100" => n11 <= "000010010110101010100000000101100011";
        when "011110101" => n11 <= "000010001010001000100000000100101010";
        when "011110110" => n11 <= "000001111101100101100000000011110110";
        when "011110111" => n11 <= "000001110001000010100000000011000111";
        when "011111000" => n11 <= "000001100100011111100000000010011101";
        when "011111001" => n11 <= "000001010111111100100000000001111000";
        when "011111010" => n11 <= "000001001011011000100000000001011000";
        when "011111011" => n11 <= "000000111110110100100000000000111101";
        when "011111100" => n11 <= "000000110010010000100000000000100111";
        when "011111101" => n11 <= "000000100101101100100000000000010110";
        when "011111110" => n11 <= "000000011001001000100000000000001001";
        when "011111111" => n11 <= "000000001100100100100000000000000010";
        when "100000000" => n11 <= "000000000000000000100000000000000000";
        when "100000001" => n11 <= "111111110011011011100000000000000010";
        when "100000010" => n11 <= "111111100110110111100000000000001001";
        when "100000011" => n11 <= "111111011010010011100000000000010110";
        when "100000100" => n11 <= "111111001101101111100000000000100111";
        when "100000101" => n11 <= "111111000001001011100000000000111101";
        when "100000110" => n11 <= "111110110100100111100000000001011000";
        when "100000111" => n11 <= "111110101000000011100000000001111000";
        when "100001000" => n11 <= "111110011011100000100000000010011101";
        when "100001001" => n11 <= "111110001110111101100000000011000111";
        when "100001010" => n11 <= "111110000010011010100000000011110110";
        when "100001011" => n11 <= "111101110101110111100000000100101010";
        when "100001100" => n11 <= "111101101001010101100000000101100011";
        when "100001101" => n11 <= "111101011100110011100000000110100000";
        when "100001110" => n11 <= "111101010000010010100000000111100011";
        when "100001111" => n11 <= "111101000011110001100000001000101010";
        when "100010000" => n11 <= "111100110111010000100000001001110111";
        when "100010001" => n11 <= "111100101010110000100000001011001000";
        when "100010010" => n11 <= "111100011110010000100000001100011110";
        when "100010011" => n11 <= "111100010001110001100000001101111001";
        when "100010100" => n11 <= "111100000101010011100000001111011001";
        when "100010101" => n11 <= "111011111000110101100000010000111110";
        when "100010110" => n11 <= "111011101100011000100000010010101000";
        when "100010111" => n11 <= "111011011111111011100000010100010111";
        when "100011000" => n11 <= "111011010011011111100000010110001010";
        when "100011001" => n11 <= "111011000111000100100000011000000011";
        when "100011010" => n11 <= "111010111010101010100000011010000000";
        when "100011011" => n11 <= "111010101110010000100000011100000010";
        when "100011100" => n11 <= "111010100001110111100000011110001001";
        when "100011101" => n11 <= "111010010101011111100000100000010101";
        when "100011110" => n11 <= "111010001001001000100000100010100110";
        when "100011111" => n11 <= "111001111100110010100000100100111100";
        when "100100000" => n11 <= "111001110000011101100000100111010110";
        when "100100001" => n11 <= "111001100100001000100000101001110101";
        when "100100010" => n11 <= "111001010111110101100000101100011001";
        when "100100011" => n11 <= "111001001011100011100000101111000010";
        when "100100100" => n11 <= "111000111111010001100000110001110000";
        when "100100101" => n11 <= "111000110011000001100000110100100011";
        when "100100110" => n11 <= "111000100110110010100000110111011010";
        when "100100111" => n11 <= "111000011010100100100000111010010111";
        when "100101000" => n11 <= "111000001110011000100000111101011000";
        when "100101001" => n11 <= "111000000010001100100001000000011101";
        when "100101010" => n11 <= "110111110110000010100001000011101000";
        when "100101011" => n11 <= "110111101001111001100001000110110111";
        when "100101100" => n11 <= "110111011101110001100001001010001011";
        when "100101101" => n11 <= "110111010001101010100001001101100100";
        when "100101110" => n11 <= "110111000101100101100001010001000010";
        when "100101111" => n11 <= "110110111001100010100001010100100100";
        when "100110000" => n11 <= "110110101101011111100001011000001011";
        when "100110001" => n11 <= "110110100001011110100001011011110111";
        when "100110010" => n11 <= "110110010101011111100001011111101000";
        when "100110011" => n11 <= "110110001001100001100001100011011101";
        when "100110100" => n11 <= "110101111101100101100001100111010111";
        when "100110101" => n11 <= "110101110001101010100001101011010110";
        when "100110110" => n11 <= "110101100101110000100001101111011001";
        when "100110111" => n11 <= "110101011001111001100001110011100001";
        when "100111000" => n11 <= "110101001110000011100001110111101101";
        when "100111001" => n11 <= "110101000010001110100001111011111111";
        when "100111010" => n11 <= "110100110110011100100010000000010101";
        when "100111011" => n11 <= "110100101010101011100010000100101111";
        when "100111100" => n11 <= "110100011110111011100010001001001110";
        when "100111101" => n11 <= "110100010011001110100010001101110010";
        when "100111110" => n11 <= "110100000111100010100010010010011010";
        when "100111111" => n11 <= "110011111011111000100010010111000111";
        when "101000000" => n11 <= "110011110000010000100010011011111001";
        when "101000001" => n11 <= "110011100100101010100010100000101111";
        when "101000010" => n11 <= "110011011001000110100010100101101001";
        when "101000011" => n11 <= "110011001101100100100010101010101001";
        when "101000100" => n11 <= "110011000010000100100010101111101100";
        when "101000101" => n11 <= "110010110110100101100010110100110100";
        when "101000110" => n11 <= "110010101011001001100010111010000001";
        when "101000111" => n11 <= "110010011111101111100010111111010010";
        when "101001000" => n11 <= "110010010100010111100011000100101000";
        when "101001001" => n11 <= "110010001001000001100011001010000010";
        when "101001010" => n11 <= "110001111101101101100011001111100000";
        when "101001011" => n11 <= "110001110010011100100011010101000011";
        when "101001100" => n11 <= "110001100111001100100011011010101011";
        when "101001101" => n11 <= "110001011011111111100011100000010111";
        when "101001110" => n11 <= "110001010000110100100011100110000111";
        when "101001111" => n11 <= "110001000101101011100011101011111011";
        when "101010000" => n11 <= "110000111010100101100011110001110100";
        when "101010001" => n11 <= "110000101111100000100011110111110010";
        when "101010010" => n11 <= "110000100100011111100011111101110011";
        when "101010011" => n11 <= "110000011001011111100100000011111001";
        when "101010100" => n11 <= "110000001110100010100100001010000011";
        when "101010101" => n11 <= "110000000011101000100100010000010010";
        when "101010110" => n11 <= "101111111000110000100100010110100101";
        when "101010111" => n11 <= "101111101101111010100100011100111100";
        when "101011000" => n11 <= "101111100011000111100100100011010111";
        when "101011001" => n11 <= "101111011000010110100100101001110111";
        when "101011010" => n11 <= "101111001101101000100100110000011011";
        when "101011011" => n11 <= "101111000010111101100100110111000011";
        when "101011100" => n11 <= "101110111000010100100100111101101111";
        when "101011101" => n11 <= "101110101101101110100101000100011111";
        when "101011110" => n11 <= "101110100011001011100101001011010100";
        when "101011111" => n11 <= "101110011000101010100101010010001100";
        when "101100000" => n11 <= "101110001110001100100101011001001001";
        when "101100001" => n11 <= "101110000011110000100101100000001010";
        when "101100010" => n11 <= "101101111001011000100101100111001111";
        when "101100011" => n11 <= "101101101111000010100101101110011000";
        when "101100100" => n11 <= "101101100100101111100101110101100101";
        when "101100101" => n11 <= "101101011010011111100101111100110110";
        when "101100110" => n11 <= "101101010000010010100110000100001011";
        when "101100111" => n11 <= "101101000110000111100110001011100100";
        when "101101000" => n11 <= "101100111100000000100110010011000001";
        when "101101001" => n11 <= "101100110001111011100110011010100011";
        when "101101010" => n11 <= "101100100111111010100110100010001000";
        when "101101011" => n11 <= "101100011101111011100110101001110001";
        when "101101100" => n11 <= "101100010100000000100110110001011101";
        when "101101101" => n11 <= "101100001010000111100110111001001110";
        when "101101110" => n11 <= "101100000000010010100111000001000011";
        when "101101111" => n11 <= "101011110110100000100111001000111011";
        when "101110000" => n11 <= "101011101100110000100111010000110111";
        when "101110001" => n11 <= "101011100011000100100111011000111000";
        when "101110010" => n11 <= "101011011001011011100111100000111011";
        when "101110011" => n11 <= "101011001111110101100111101001000011";
        when "101110100" => n11 <= "101011000110010011100111110001001111";
        when "101110101" => n11 <= "101010111100110011100111111001011110";
        when "101110110" => n11 <= "101010110011010111101000000001110001";
        when "101110111" => n11 <= "101010101001111110101000001010000111";
        when "101111000" => n11 <= "101010100000101001101000010010100010";
        when "101111001" => n11 <= "101010010111010111101000011010111111";
        when "101111010" => n11 <= "101010001110001000101000100011100001";
        when "101111011" => n11 <= "101010000100111100101000101100000110";
        when "101111100" => n11 <= "101001111011110100101000110100101111";
        when "101111101" => n11 <= "101001110010101111101000111101011011";
        when "101111110" => n11 <= "101001101001101110101001000110001011";
        when "101111111" => n11 <= "101001100000110000101001001110111111";
        when "110000000" => n11 <= "101001010111110110101001010111110110";
        when "110000001" => n11 <= "101001001110111111101001100000110000";
        when "110000010" => n11 <= "101001000110001011101001101001101110";
        when "110000011" => n11 <= "101000111101011011101001110010101111";
        when "110000100" => n11 <= "101000110100101111101001111011110100";
        when "110000101" => n11 <= "101000101100000110101010000100111100";
        when "110000110" => n11 <= "101000100011100001101010001110001000";
        when "110000111" => n11 <= "101000011010111111101010010111010111";
        when "110001000" => n11 <= "101000010010100010101010100000101001";
        when "110001001" => n11 <= "101000001010000111101010101001111110";
        when "110001010" => n11 <= "101000000001110001101010110011010111";
        when "110001011" => n11 <= "100111111001011110101010111100110011";
        when "110001100" => n11 <= "100111110001001111101011000110010011";
        when "110001101" => n11 <= "100111101001000011101011001111110101";
        when "110001110" => n11 <= "100111100000111011101011011001011011";
        when "110001111" => n11 <= "100111011000111000101011100011000100";
        when "110010000" => n11 <= "100111010000110111101011101100110000";
        when "110010001" => n11 <= "100111001000111011101011110110100000";
        when "110010010" => n11 <= "100111000001000011101100000000010010";
        when "110010011" => n11 <= "100110111001001110101100001010000111";
        when "110010100" => n11 <= "100110110001011101101100010100000000";
        when "110010101" => n11 <= "100110101001110001101100011101111011";
        when "110010110" => n11 <= "100110100010001000101100100111111010";
        when "110010111" => n11 <= "100110011010100011101100110001111011";
        when "110011000" => n11 <= "100110010011000001101100111100000000";
        when "110011001" => n11 <= "100110001011100100101101000110000111";
        when "110011010" => n11 <= "100110000100001011101101010000010010";
        when "110011011" => n11 <= "100101111100110110101101011010011111";
        when "110011100" => n11 <= "100101110101100101101101100100101111";
        when "110011101" => n11 <= "100101101110011000101101101111000010";
        when "110011110" => n11 <= "100101100111001111101101111001011000";
        when "110011111" => n11 <= "100101100000001010101110000011110000";
        when "110100000" => n11 <= "100101011001001001101110001110001100";
        when "110100001" => n11 <= "100101010010001100101110011000101010";
        when "110100010" => n11 <= "100101001011010100101110100011001011";
        when "110100011" => n11 <= "100101000100011111101110101101101110";
        when "110100100" => n11 <= "100100111101101111101110111000010100";
        when "110100101" => n11 <= "100100110111000011101111000010111101";
        when "110100110" => n11 <= "100100110000011011101111001101101000";
        when "110100111" => n11 <= "100100101001110111101111011000010110";
        when "110101000" => n11 <= "100100100011010111101111100011000111";
        when "110101001" => n11 <= "100100011100111100101111101101111010";
        when "110101010" => n11 <= "100100010110100101101111111000110000";
        when "110101011" => n11 <= "100100010000010010110000000011101000";
        when "110101100" => n11 <= "100100001010000011110000001110100010";
        when "110101101" => n11 <= "100100000011111001110000011001011111";
        when "110101110" => n11 <= "100011111101110011110000100100011111";
        when "110101111" => n11 <= "100011110111110010110000101111100000";
        when "110110000" => n11 <= "100011110001110100110000111010100101";
        when "110110001" => n11 <= "100011101011111011110001000101101011";
        when "110110010" => n11 <= "100011100110000111110001010000110100";
        when "110110011" => n11 <= "100011100000010111110001011011111111";
        when "110110100" => n11 <= "100011011010101011110001100111001100";
        when "110110101" => n11 <= "100011010101000011110001110010011100";
        when "110110110" => n11 <= "100011001111100000110001111101101101";
        when "110110111" => n11 <= "100011001010000010110010001001000001";
        when "110111000" => n11 <= "100011000100101000110010010100010111";
        when "110111001" => n11 <= "100010111111010010110010011111101111";
        when "110111010" => n11 <= "100010111010000001110010101011001001";
        when "110111011" => n11 <= "100010110100110100110010110110100101";
        when "110111100" => n11 <= "100010101111101100110011000010000100";
        when "110111101" => n11 <= "100010101010101001110011001101100100";
        when "110111110" => n11 <= "100010100101101001110011011001000110";
        when "110111111" => n11 <= "100010100000101111110011100100101010";
        when "111000000" => n11 <= "100010011011111001110011110000010000";
        when "111000001" => n11 <= "100010010111000111110011111011111000";
        when "111000010" => n11 <= "100010010010011010110100000111100010";
        when "111000011" => n11 <= "100010001101110010110100010011001110";
        when "111000100" => n11 <= "100010001001001110110100011110111011";
        when "111000101" => n11 <= "100010000100101111110100101010101011";
        when "111000110" => n11 <= "100010000000010101110100110110011100";
        when "111000111" => n11 <= "100001111011111111110101000010001110";
        when "111001000" => n11 <= "100001110111101101110101001110000011";
        when "111001001" => n11 <= "100001110011100001110101011001111001";
        when "111001010" => n11 <= "100001101111011001110101100101110000";
        when "111001011" => n11 <= "100001101011010110110101110001101010";
        when "111001100" => n11 <= "100001100111010111110101111101100101";
        when "111001101" => n11 <= "100001100011011101110110001001100001";
        when "111001110" => n11 <= "100001011111101000110110010101011111";
        when "111001111" => n11 <= "100001011011110111110110100001011110";
        when "111010000" => n11 <= "100001011000001011110110101101011111";
        when "111010001" => n11 <= "100001010100100100110110111001100010";
        when "111010010" => n11 <= "100001010001000010110111000101100101";
        when "111010011" => n11 <= "100001001101100100110111010001101010";
        when "111010100" => n11 <= "100001001010001011110111011101110001";
        when "111010101" => n11 <= "100001000110110111110111101001111001";
        when "111010110" => n11 <= "100001000011101000110111110110000010";
        when "111010111" => n11 <= "100001000000011101111000000010001100";
        when "111011000" => n11 <= "100000111101011000111000001110011000";
        when "111011001" => n11 <= "100000111010010111111000011010100100";
        when "111011010" => n11 <= "100000110111011010111000100110110010";
        when "111011011" => n11 <= "100000110100100011111000110011000001";
        when "111011100" => n11 <= "100000110001110000111000111111010001";
        when "111011101" => n11 <= "100000101111000010111001001011100011";
        when "111011110" => n11 <= "100000101100011001111001010111110101";
        when "111011111" => n11 <= "100000101001110101111001100100001000";
        when "111100000" => n11 <= "100000100111010110111001110000011101";
        when "111100001" => n11 <= "100000100100111100111001111100110010";
        when "111100010" => n11 <= "100000100010100110111010001001001000";
        when "111100011" => n11 <= "100000100000010101111010010101011111";
        when "111100100" => n11 <= "100000011110001001111010100001110111";
        when "111100101" => n11 <= "100000011100000010111010101110010000";
        when "111100110" => n11 <= "100000011010000000111010111010101010";
        when "111100111" => n11 <= "100000011000000011111011000111000100";
        when "111101000" => n11 <= "100000010110001010111011010011011111";
        when "111101001" => n11 <= "100000010100010111111011011111111011";
        when "111101010" => n11 <= "100000010010101000111011101100011000";
        when "111101011" => n11 <= "100000010000111110111011111000110101";
        when "111101100" => n11 <= "100000001111011001111100000101010011";
        when "111101101" => n11 <= "100000001101111001111100010001110001";
        when "111101110" => n11 <= "100000001100011110111100011110010000";
        when "111101111" => n11 <= "100000001011001000111100101010110000";
        when "111110000" => n11 <= "100000001001110111111100110111010000";
        when "111110001" => n11 <= "100000001000101010111101000011110001";
        when "111110010" => n11 <= "100000000111100011111101010000010010";
        when "111110011" => n11 <= "100000000110100000111101011100110011";
        when "111110100" => n11 <= "100000000101100011111101101001010101";
        when "111110101" => n11 <= "100000000100101010111101110101110111";
        when "111110110" => n11 <= "100000000011110110111110000010011010";
        when "111110111" => n11 <= "100000000011000111111110001110111101";
        when "111111000" => n11 <= "100000000010011101111110011011100000";
        when "111111001" => n11 <= "100000000001111000111110101000000011";
        when "111111010" => n11 <= "100000000001011000111110110100100111";
        when "111111011" => n11 <= "100000000000111101111111000001001011";
        when "111111100" => n11 <= "100000000000100111111111001101101111";
        when "111111101" => n11 <= "100000000000010110111111011010010011";
        when "111111110" => n11 <= "100000000000001001111111100110110111";
        when "111111111" => n11 <= "100000000000000010111111110011011011";
        when others => n11 <= "XXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX";
      end case;
    end if;
  end if;
end process;
n12 <= n11(35 downto 35) &
  n11(34 downto 34) &
  n11(33 downto 33) &
  n11(32 downto 32) &
  n11(31 downto 31) &
  n11(30 downto 30) &
  n11(29 downto 29) &
  n11(28 downto 28) &
  n11(27 downto 27) &
  n11(26 downto 26) &
  n11(25 downto 25) &
  n11(24 downto 24) &
  n11(23 downto 23) &
  n11(22 downto 22) &
  n11(21 downto 21) &
  n11(20 downto 20) &
  n11(19 downto 19) &
  n11(18 downto 18);
n13 <= n11(17 downto 17) &
  n11(16 downto 16) &
  n11(15 downto 15) &
  n11(14 downto 14) &
  n11(13 downto 13) &
  n11(12 downto 12) &
  n11(11 downto 11) &
  n11(10 downto 10) &
  n11(9 downto 9) &
  n11(8 downto 8) &
  n11(7 downto 7) &
  n11(6 downto 6) &
  n11(5 downto 5) &
  n11(4 downto 4) &
  n11(3 downto 3) &
  n11(2 downto 2) &
  n11(1 downto 1) &
  n11(0 downto 0);
n14 <= unsigned(signed(n5) * signed(n12));
n15 <= n14(34 downto 34) &
  n14(33 downto 33) &
  n14(32 downto 32) &
  n14(31 downto 31) &
  n14(30 downto 30) &
  n14(29 downto 29) &
  n14(28 downto 28) &
  n14(27 downto 27) &
  n14(26 downto 26) &
  n14(25 downto 25) &
  n14(24 downto 24) &
  n14(23 downto 23) &
  n14(22 downto 22) &
  n14(21 downto 21) &
  n14(20 downto 20) &
  n14(19 downto 19) &
  n14(18 downto 18) &
  n14(17 downto 17);
process (clock_c) begin
  if rising_edge(clock_c) then
    if i5 = "1" then
      n16 <= "000000000000000000";
    elsif i4 = "1" then
      n16 <= n15;
    end if;
  end if;
end process;
n17 <= unsigned(signed(n6) * signed(n13));
n18 <= n17(34 downto 34) &
  n17(33 downto 33) &
  n17(32 downto 32) &
  n17(31 downto 31) &
  n17(30 downto 30) &
  n17(29 downto 29) &
  n17(28 downto 28) &
  n17(27 downto 27) &
  n17(26 downto 26) &
  n17(25 downto 25) &
  n17(24 downto 24) &
  n17(23 downto 23) &
  n17(22 downto 22) &
  n17(21 downto 21) &
  n17(20 downto 20) &
  n17(19 downto 19) &
  n17(18 downto 18) &
  n17(17 downto 17);
process (clock_c) begin
  if rising_edge(clock_c) then
    if i5 = "1" then
      n19 <= "000000000000000000";
    elsif i4 = "1" then
      n19 <= n18;
    end if;
  end if;
end process;
n20 <= n16 - n19;
process (clock_c) begin
  if rising_edge(clock_c) then
    if i5 = "1" then
      n21 <= "000000000000000000";
    elsif i4 = "1" then
      n21 <= n20;
    end if;
  end if;
end process;
n22 <= unsigned(signed(n5) * signed(n13));
n23 <= n22(34 downto 34) &
  n22(33 downto 33) &
  n22(32 downto 32) &
  n22(31 downto 31) &
  n22(30 downto 30) &
  n22(29 downto 29) &
  n22(28 downto 28) &
  n22(27 downto 27) &
  n22(26 downto 26) &
  n22(25 downto 25) &
  n22(24 downto 24) &
  n22(23 downto 23) &
  n22(22 downto 22) &
  n22(21 downto 21) &
  n22(20 downto 20) &
  n22(19 downto 19) &
  n22(18 downto 18) &
  n22(17 downto 17);
process (clock_c) begin
  if rising_edge(clock_c) then
    if i5 = "1" then
      n24 <= "000000000000000000";
    elsif i4 = "1" then
      n24 <= n23;
    end if;
  end if;
end process;
n25 <= unsigned(signed(n6) * signed(n12));
n26 <= n25(34 downto 34) &
  n25(33 downto 33) &
  n25(32 downto 32) &
  n25(31 downto 31) &
  n25(30 downto 30) &
  n25(29 downto 29) &
  n25(28 downto 28) &
  n25(27 downto 27) &
  n25(26 downto 26) &
  n25(25 downto 25) &
  n25(24 downto 24) &
  n25(23 downto 23) &
  n25(22 downto 22) &
  n25(21 downto 21) &
  n25(20 downto 20) &
  n25(19 downto 19) &
  n25(18 downto 18) &
  n25(17 downto 17);
process (clock_c) begin
  if rising_edge(clock_c) then
    if i5 = "1" then
      n27 <= "000000000000000000";
    elsif i4 = "1" then
      n27 <= n26;
    end if;
  end if;
end process;
n28 <= n24 + n27;
process (clock_c) begin
  if rising_edge(clock_c) then
    if i5 = "1" then
      n29 <= "000000000000000000";
    elsif i4 = "1" then
      n29 <= n28;
    end if;
  end if;
end process;
n30 <= n8 + n21;
n31 <= n10 + n29;
n32 <= n30 & n31;
process (clock_c) begin
  if rising_edge(clock_c) then
    if i5 = "1" then
      n33 <= "000000000000000000000000000000000000";
    elsif i4 = "1" then
      n33 <= n32;
    end if;
  end if;
end process;
n34 <= n8 - n21;
n35 <= n10 - n29;
n36 <= n34 & n35;
process (clock_c) begin
  if rising_edge(clock_c) then
    if i5 = "1" then
      n37 <= "000000000000000000000000000000000000";
    elsif i4 = "1" then
      n37 <= n36;
    end if;
  end if;
end process;
o2 <= n37;
o1 <= n33;
end architecture rtl;

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
entity cf_fft_4096_18_21 is
port (
clock_c : in std_logic;
i1 : in  unsigned(0 downto 0);
i2 : in  unsigned(35 downto 0);
i3 : in  unsigned(35 downto 0);
i4 : in  unsigned(0 downto 0);
i5 : in  unsigned(0 downto 0);
o1 : out unsigned(0 downto 0);
o2 : out unsigned(35 downto 0);
o3 : out unsigned(35 downto 0));
end entity cf_fft_4096_18_21;
architecture rtl of cf_fft_4096_18_21 is
signal n1 : unsigned(8 downto 0);
signal n2 : unsigned(71 downto 0);
signal n3 : unsigned(0 downto 0) := "0";
signal n4 : unsigned(0 downto 0) := "0";
signal n5 : unsigned(0 downto 0) := "0";
signal n6 : unsigned(0 downto 0) := "0";
signal n7 : unsigned(9 downto 0);
signal n8 : unsigned(9 downto 0) := "0000000000";
signal n9 : unsigned(9 downto 0) := "0000000000";
signal n10 : unsigned(9 downto 0) := "0000000000";
signal n11 : unsigned(9 downto 0) := "0000000000";
signal n12 : unsigned(0 downto 0);
signal n13 : unsigned(0 downto 0) := "0";
signal n14 : unsigned(0 downto 0) := "0";
signal n15 : unsigned(0 downto 0) := "0";
signal n16 : unsigned(0 downto 0) := "0";
signal n17 : unsigned(0 downto 0);
signal n18 : unsigned(1 downto 0);
signal n19 : unsigned(35 downto 0);
signal n20 : unsigned(35 downto 0);
signal n21 : unsigned(35 downto 0);
signal n22 : unsigned(35 downto 0);
signal n23 : unsigned(35 downto 0);
signal n24 : unsigned(35 downto 0);
signal s25_1 : unsigned(35 downto 0);
signal s25_2 : unsigned(35 downto 0);
signal s26_1 : unsigned(0 downto 0);
signal s27_1 : unsigned(71 downto 0);
signal s28_1 : unsigned(0 downto 0);
signal s28_2 : unsigned(0 downto 0);
signal s28_3 : unsigned(71 downto 0);
signal s29_1 : unsigned(10 downto 0);
signal s29_2 : unsigned(0 downto 0);
component cf_fft_4096_18_22 is
port (
clock_c : in std_logic;
i1 : in  unsigned(35 downto 0);
i2 : in  unsigned(35 downto 0);
i3 : in  unsigned(8 downto 0);
i4 : in  unsigned(0 downto 0);
i5 : in  unsigned(0 downto 0);
o1 : out unsigned(35 downto 0);
o2 : out unsigned(35 downto 0));
end component cf_fft_4096_18_22;
component cf_fft_4096_18_37 is
port (
clock_c : in std_logic;
i1 : in  unsigned(1 downto 0);
i2 : in  unsigned(0 downto 0);
i3 : in  unsigned(0 downto 0);
o1 : out unsigned(0 downto 0));
end component cf_fft_4096_18_37;
component cf_fft_4096_18_33 is
port (
clock_c : in std_logic;
i1 : in  unsigned(71 downto 0);
i2 : in  unsigned(0 downto 0);
i3 : in  unsigned(9 downto 0);
i4 : in  unsigned(0 downto 0);
i5 : in  unsigned(0 downto 0);
i6 : in  unsigned(0 downto 0);
o1 : out unsigned(71 downto 0));
end component cf_fft_4096_18_33;
component cf_fft_4096_18_32 is
port (
clock_c : in std_logic;
i1 : in  unsigned(71 downto 0);
i2 : in  unsigned(0 downto 0);
i3 : in  unsigned(9 downto 0);
i4 : in  unsigned(0 downto 0);
i5 : in  unsigned(0 downto 0);
i6 : in  unsigned(0 downto 0);
o1 : out unsigned(0 downto 0);
o2 : out unsigned(0 downto 0);
o3 : out unsigned(71 downto 0));
end component cf_fft_4096_18_32;
component cf_fft_4096_18_28 is
port (
clock_c : in std_logic;
i1 : in  unsigned(0 downto 0);
i2 : in  unsigned(0 downto 0);
i3 : in  unsigned(0 downto 0);
o1 : out unsigned(10 downto 0);
o2 : out unsigned(0 downto 0));
end component cf_fft_4096_18_28;
begin
n1 <= s29_1(10 downto 10) &
  s29_1(9 downto 9) &
  s29_1(8 downto 8) &
  s29_1(7 downto 7) &
  s29_1(6 downto 6) &
  s29_1(5 downto 5) &
  s29_1(4 downto 4) &
  s29_1(3 downto 3) &
  s29_1(2 downto 2);
n2 <= s25_1 & s25_2;
process (clock_c) begin
  if rising_edge(clock_c) then
    if i5 = "1" then
      n3 <= "0";
    elsif i4 = "1" then
      n3 <= s29_2;
    end if;
  end if;
end process;
process (clock_c) begin
  if rising_edge(clock_c) then
    if i5 = "1" then
      n4 <= "0";
    elsif i4 = "1" then
      n4 <= n3;
    end if;
  end if;
end process;
process (clock_c) begin
  if rising_edge(clock_c) then
    if i5 = "1" then
      n5 <= "0";
    elsif i4 = "1" then
      n5 <= n4;
    end if;
  end if;
end process;
process (clock_c) begin
  if rising_edge(clock_c) then
    if i5 = "1" then
      n6 <= "0";
    elsif i4 = "1" then
      n6 <= n5;
    end if;
  end if;
end process;
n7 <= s29_1(10 downto 10) &
  s29_1(9 downto 9) &
  s29_1(8 downto 8) &
  s29_1(7 downto 7) &
  s29_1(6 downto 6) &
  s29_1(5 downto 5) &
  s29_1(4 downto 4) &
  s29_1(3 downto 3) &
  s29_1(2 downto 2) &
  s29_1(1 downto 1);
process (clock_c) begin
  if rising_edge(clock_c) then
    if i5 = "1" then
      n8 <= "0000000000";
    elsif i4 = "1" then
      n8 <= n7;
    end if;
  end if;
end process;
process (clock_c) begin
  if rising_edge(clock_c) then
    if i5 = "1" then
      n9 <= "0000000000";
    elsif i4 = "1" then
      n9 <= n8;
    end if;
  end if;
end process;
process (clock_c) begin
  if rising_edge(clock_c) then
    if i5 = "1" then
      n10 <= "0000000000";
    elsif i4 = "1" then
      n10 <= n9;
    end if;
  end if;
end process;
process (clock_c) begin
  if rising_edge(clock_c) then
    if i5 = "1" then
      n11 <= "0000000000";
    elsif i4 = "1" then
      n11 <= n10;
    end if;
  end if;
end process;
n12 <= s29_1(0 downto 0);
process (clock_c) begin
  if rising_edge(clock_c) then
    if i5 = "1" then
      n13 <= "0";
    elsif i4 = "1" then
      n13 <= n12;
    end if;
  end if;
end process;
process (clock_c) begin
  if rising_edge(clock_c) then
    if i5 = "1" then
      n14 <= "0";
    elsif i4 = "1" then
      n14 <= n13;
    end if;
  end if;
end process;
process (clock_c) begin
  if rising_edge(clock_c) then
    if i5 = "1" then
      n15 <= "0";
    elsif i4 = "1" then
      n15 <= n14;
    end if;
  end if;
end process;
process (clock_c) begin
  if rising_edge(clock_c) then
    if i5 = "1" then
      n16 <= "0";
    elsif i4 = "1" then
      n16 <= n15;
    end if;
  end if;
end process;
n17 <= not n16;
n18 <= s28_2 & s28_1;
n19 <= s28_3(71 downto 71) &
  s28_3(70 downto 70) &
  s28_3(69 downto 69) &
  s28_3(68 downto 68) &
  s28_3(67 downto 67) &
  s28_3(66 downto 66) &
  s28_3(65 downto 65) &
  s28_3(64 downto 64) &
  s28_3(63 downto 63) &
  s28_3(62 downto 62) &
  s28_3(61 downto 61) &
  s28_3(60 downto 60) &
  s28_3(59 downto 59) &
  s28_3(58 downto 58) &
  s28_3(57 downto 57) &
  s28_3(56 downto 56) &
  s28_3(55 downto 55) &
  s28_3(54 downto 54) &
  s28_3(53 downto 53) &
  s28_3(52 downto 52) &
  s28_3(51 downto 51) &
  s28_3(50 downto 50) &
  s28_3(49 downto 49) &
  s28_3(48 downto 48) &
  s28_3(47 downto 47) &
  s28_3(46 downto 46) &
  s28_3(45 downto 45) &
  s28_3(44 downto 44) &
  s28_3(43 downto 43) &
  s28_3(42 downto 42) &
  s28_3(41 downto 41) &
  s28_3(40 downto 40) &
  s28_3(39 downto 39) &
  s28_3(38 downto 38) &
  s28_3(37 downto 37) &
  s28_3(36 downto 36);
n20 <= s28_3(35 downto 35) &
  s28_3(34 downto 34) &
  s28_3(33 downto 33) &
  s28_3(32 downto 32) &
  s28_3(31 downto 31) &
  s28_3(30 downto 30) &
  s28_3(29 downto 29) &
  s28_3(28 downto 28) &
  s28_3(27 downto 27) &
  s28_3(26 downto 26) &
  s28_3(25 downto 25) &
  s28_3(24 downto 24) &
  s28_3(23 downto 23) &
  s28_3(22 downto 22) &
  s28_3(21 downto 21) &
  s28_3(20 downto 20) &
  s28_3(19 downto 19) &
  s28_3(18 downto 18) &
  s28_3(17 downto 17) &
  s28_3(16 downto 16) &
  s28_3(15 downto 15) &
  s28_3(14 downto 14) &
  s28_3(13 downto 13) &
  s28_3(12 downto 12) &
  s28_3(11 downto 11) &
  s28_3(10 downto 10) &
  s28_3(9 downto 9) &
  s28_3(8 downto 8) &
  s28_3(7 downto 7) &
  s28_3(6 downto 6) &
  s28_3(5 downto 5) &
  s28_3(4 downto 4) &
  s28_3(3 downto 3) &
  s28_3(2 downto 2) &
  s28_3(1 downto 1) &
  s28_3(0 downto 0);
n21 <= s27_1(71 downto 71) &
  s27_1(70 downto 70) &
  s27_1(69 downto 69) &
  s27_1(68 downto 68) &
  s27_1(67 downto 67) &
  s27_1(66 downto 66) &
  s27_1(65 downto 65) &
  s27_1(64 downto 64) &
  s27_1(63 downto 63) &
  s27_1(62 downto 62) &
  s27_1(61 downto 61) &
  s27_1(60 downto 60) &
  s27_1(59 downto 59) &
  s27_1(58 downto 58) &
  s27_1(57 downto 57) &
  s27_1(56 downto 56) &
  s27_1(55 downto 55) &
  s27_1(54 downto 54) &
  s27_1(53 downto 53) &
  s27_1(52 downto 52) &
  s27_1(51 downto 51) &
  s27_1(50 downto 50) &
  s27_1(49 downto 49) &
  s27_1(48 downto 48) &
  s27_1(47 downto 47) &
  s27_1(46 downto 46) &
  s27_1(45 downto 45) &
  s27_1(44 downto 44) &
  s27_1(43 downto 43) &
  s27_1(42 downto 42) &
  s27_1(41 downto 41) &
  s27_1(40 downto 40) &
  s27_1(39 downto 39) &
  s27_1(38 downto 38) &
  s27_1(37 downto 37) &
  s27_1(36 downto 36);
n22 <= s27_1(35 downto 35) &
  s27_1(34 downto 34) &
  s27_1(33 downto 33) &
  s27_1(32 downto 32) &
  s27_1(31 downto 31) &
  s27_1(30 downto 30) &
  s27_1(29 downto 29) &
  s27_1(28 downto 28) &
  s27_1(27 downto 27) &
  s27_1(26 downto 26) &
  s27_1(25 downto 25) &
  s27_1(24 downto 24) &
  s27_1(23 downto 23) &
  s27_1(22 downto 22) &
  s27_1(21 downto 21) &
  s27_1(20 downto 20) &
  s27_1(19 downto 19) &
  s27_1(18 downto 18) &
  s27_1(17 downto 17) &
  s27_1(16 downto 16) &
  s27_1(15 downto 15) &
  s27_1(14 downto 14) &
  s27_1(13 downto 13) &
  s27_1(12 downto 12) &
  s27_1(11 downto 11) &
  s27_1(10 downto 10) &
  s27_1(9 downto 9) &
  s27_1(8 downto 8) &
  s27_1(7 downto 7) &
  s27_1(6 downto 6) &
  s27_1(5 downto 5) &
  s27_1(4 downto 4) &
  s27_1(3 downto 3) &
  s27_1(2 downto 2) &
  s27_1(1 downto 1) &
  s27_1(0 downto 0);
n23 <= n20 when s26_1 = "1" else n19;
n24 <= n22 when s26_1 = "1" else n21;
s25 : cf_fft_4096_18_22 port map (clock_c, i2, i3, n1, i4, i5, s25_1, s25_2);
s26 : cf_fft_4096_18_37 port map (clock_c, n18, i4, i5, s26_1);
s27 : cf_fft_4096_18_33 port map (clock_c, n2, n6, n11, n16, i4, i5, s27_1);
s28 : cf_fft_4096_18_32 port map (clock_c, n2, n6, n11, n17, i4, i5, s28_1, s28_2, s28_3);
s29 : cf_fft_4096_18_28 port map (clock_c, i1, i4, i5, s29_1, s29_2);
o3 <= n24;
o2 <= n23;
o1 <= s28_1;
end architecture rtl;

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
entity cf_fft_4096_18_20 is
port (
clock_c : in std_logic;
i1 : in  unsigned(35 downto 0);
i2 : in  unsigned(35 downto 0);
i3 : in  unsigned(7 downto 0);
i4 : in  unsigned(0 downto 0);
i5 : in  unsigned(0 downto 0);
o1 : out unsigned(35 downto 0);
o2 : out unsigned(35 downto 0));
end entity cf_fft_4096_18_20;
architecture rtl of cf_fft_4096_18_20 is
signal n1 : unsigned(35 downto 0) := "000000000000000000000000000000000000";
signal n2 : unsigned(17 downto 0);
signal n3 : unsigned(17 downto 0);
signal n4 : unsigned(35 downto 0) := "000000000000000000000000000000000000";
signal n5 : unsigned(17 downto 0);
signal n6 : unsigned(17 downto 0);
signal n7 : unsigned(17 downto 0) := "000000000000000000";
signal n8 : unsigned(17 downto 0) := "000000000000000000";
signal n9 : unsigned(17 downto 0) := "000000000000000000";
signal n10 : unsigned(17 downto 0) := "000000000000000000";
signal n11 : unsigned(35 downto 0) := "000000000000000000000000000000000000";
signal n12 : unsigned(17 downto 0);
signal n13 : unsigned(17 downto 0);
signal n14 : unsigned(35 downto 0);
signal n15 : unsigned(17 downto 0);
signal n16 : unsigned(17 downto 0) := "000000000000000000";
signal n17 : unsigned(35 downto 0);
signal n18 : unsigned(17 downto 0);
signal n19 : unsigned(17 downto 0) := "000000000000000000";
signal n20 : unsigned(17 downto 0);
signal n21 : unsigned(17 downto 0) := "000000000000000000";
signal n22 : unsigned(35 downto 0);
signal n23 : unsigned(17 downto 0);
signal n24 : unsigned(17 downto 0) := "000000000000000000";
signal n25 : unsigned(35 downto 0);
signal n26 : unsigned(17 downto 0);
signal n27 : unsigned(17 downto 0) := "000000000000000000";
signal n28 : unsigned(17 downto 0);
signal n29 : unsigned(17 downto 0) := "000000000000000000";
signal n30 : unsigned(17 downto 0);
signal n31 : unsigned(17 downto 0);
signal n32 : unsigned(35 downto 0);
signal n33 : unsigned(35 downto 0) := "000000000000000000000000000000000000";
signal n34 : unsigned(17 downto 0);
signal n35 : unsigned(17 downto 0);
signal n36 : unsigned(35 downto 0);
signal n37 : unsigned(35 downto 0) := "000000000000000000000000000000000000";
begin
process (clock_c) begin
  if rising_edge(clock_c) then
    if i5 = "1" then
      n1 <= "000000000000000000000000000000000000";
    elsif i4 = "1" then
      n1 <= i1;
    end if;
  end if;
end process;
n2 <= n1(35 downto 35) &
  n1(34 downto 34) &
  n1(33 downto 33) &
  n1(32 downto 32) &
  n1(31 downto 31) &
  n1(30 downto 30) &
  n1(29 downto 29) &
  n1(28 downto 28) &
  n1(27 downto 27) &
  n1(26 downto 26) &
  n1(25 downto 25) &
  n1(24 downto 24) &
  n1(23 downto 23) &
  n1(22 downto 22) &
  n1(21 downto 21) &
  n1(20 downto 20) &
  n1(19 downto 19) &
  n1(18 downto 18);
n3 <= n1(17 downto 17) &
  n1(16 downto 16) &
  n1(15 downto 15) &
  n1(14 downto 14) &
  n1(13 downto 13) &
  n1(12 downto 12) &
  n1(11 downto 11) &
  n1(10 downto 10) &
  n1(9 downto 9) &
  n1(8 downto 8) &
  n1(7 downto 7) &
  n1(6 downto 6) &
  n1(5 downto 5) &
  n1(4 downto 4) &
  n1(3 downto 3) &
  n1(2 downto 2) &
  n1(1 downto 1) &
  n1(0 downto 0);
process (clock_c) begin
  if rising_edge(clock_c) then
    if i5 = "1" then
      n4 <= "000000000000000000000000000000000000";
    elsif i4 = "1" then
      n4 <= i2;
    end if;
  end if;
end process;
n5 <= n4(35 downto 35) &
  n4(34 downto 34) &
  n4(33 downto 33) &
  n4(32 downto 32) &
  n4(31 downto 31) &
  n4(30 downto 30) &
  n4(29 downto 29) &
  n4(28 downto 28) &
  n4(27 downto 27) &
  n4(26 downto 26) &
  n4(25 downto 25) &
  n4(24 downto 24) &
  n4(23 downto 23) &
  n4(22 downto 22) &
  n4(21 downto 21) &
  n4(20 downto 20) &
  n4(19 downto 19) &
  n4(18 downto 18);
n6 <= n4(17 downto 17) &
  n4(16 downto 16) &
  n4(15 downto 15) &
  n4(14 downto 14) &
  n4(13 downto 13) &
  n4(12 downto 12) &
  n4(11 downto 11) &
  n4(10 downto 10) &
  n4(9 downto 9) &
  n4(8 downto 8) &
  n4(7 downto 7) &
  n4(6 downto 6) &
  n4(5 downto 5) &
  n4(4 downto 4) &
  n4(3 downto 3) &
  n4(2 downto 2) &
  n4(1 downto 1) &
  n4(0 downto 0);
process (clock_c) begin
  if rising_edge(clock_c) then
    if i5 = "1" then
      n7 <= "000000000000000000";
    elsif i4 = "1" then
      n7 <= n2;
    end if;
  end if;
end process;
process (clock_c) begin
  if rising_edge(clock_c) then
    if i5 = "1" then
      n8 <= "000000000000000000";
    elsif i4 = "1" then
      n8 <= n7;
    end if;
  end if;
end process;
process (clock_c) begin
  if rising_edge(clock_c) then
    if i5 = "1" then
      n9 <= "000000000000000000";
    elsif i4 = "1" then
      n9 <= n3;
    end if;
  end if;
end process;
process (clock_c) begin
  if rising_edge(clock_c) then
    if i5 = "1" then
      n10 <= "000000000000000000";
    elsif i4 = "1" then
      n10 <= n9;
    end if;
  end if;
end process;
process (clock_c) begin
  if rising_edge(clock_c) then 
    if i4 = "1" then
      case i3 is
        when "00000000" => n11 <= "011111111111111111000000000000000000";
        when "00000001" => n11 <= "011111111111110110111111100110110111";
        when "00000010" => n11 <= "011111111111011000111111001101101111";
        when "00000011" => n11 <= "011111111110100111111110110100100111";
        when "00000100" => n11 <= "011111111101100010111110011011100000";
        when "00000101" => n11 <= "011111111100001001111110000010011010";
        when "00000110" => n11 <= "011111111010011100111101101001010101";
        when "00000111" => n11 <= "011111111000011100111101010000010010";
        when "00001000" => n11 <= "011111110110001000111100110111010000";
        when "00001001" => n11 <= "011111110011100001111100011110010000";
        when "00001010" => n11 <= "011111110000100110111100000101010011";
        when "00001011" => n11 <= "011111101101010111111011101100011000";
        when "00001100" => n11 <= "011111101001110101111011010011011111";
        when "00001101" => n11 <= "011111100101111111111010111010101010";
        when "00001110" => n11 <= "011111100001110110111010100001110111";
        when "00001111" => n11 <= "011111011101011001111010001001001000";
        when "00010000" => n11 <= "011111011000101001111001110000011101";
        when "00010001" => n11 <= "011111010011100110111001010111110101";
        when "00010010" => n11 <= "011111001110001111111000111111010001";
        when "00010011" => n11 <= "011111001000100101111000100110110010";
        when "00010100" => n11 <= "011111000010100111111000001110011000";
        when "00010101" => n11 <= "011110111100010111110111110110000010";
        when "00010110" => n11 <= "011110110101110100110111011101110001";
        when "00010111" => n11 <= "011110101110111101110111000101100101";
        when "00011000" => n11 <= "011110100111110100110110101101011111";
        when "00011001" => n11 <= "011110100000010111110110010101011111";
        when "00011010" => n11 <= "011110011000101000110101111101100101";
        when "00011011" => n11 <= "011110010000100110110101100101110000";
        when "00011100" => n11 <= "011110001000010010110101001110000011";
        when "00011101" => n11 <= "011101111111101010110100110110011100";
        when "00011110" => n11 <= "011101110110110001110100011110111011";
        when "00011111" => n11 <= "011101101101100101110100000111100010";
        when "00100000" => n11 <= "011101100100000110110011110000010000";
        when "00100001" => n11 <= "011101011010010110110011011001000110";
        when "00100010" => n11 <= "011101010000010011110011000010000100";
        when "00100011" => n11 <= "011101000101111110110010101011001001";
        when "00100100" => n11 <= "011100111011010111110010010100010111";
        when "00100101" => n11 <= "011100110000011111110001111101101101";
        when "00100110" => n11 <= "011100100101010100110001100111001100";
        when "00100111" => n11 <= "011100011001111000110001010000110100";
        when "00101000" => n11 <= "011100001110001011110000111010100101";
        when "00101001" => n11 <= "011100000010001100110000100100011111";
        when "00101010" => n11 <= "011011110101111100110000001110100010";
        when "00101011" => n11 <= "011011101001011010101111111000110000";
        when "00101100" => n11 <= "011011011100101000101111100011000111";
        when "00101101" => n11 <= "011011001111100100101111001101101000";
        when "00101110" => n11 <= "011011000010010000101110111000010100";
        when "00101111" => n11 <= "011010110100101011101110100011001011";
        when "00110000" => n11 <= "011010100110110110101110001110001100";
        when "00110001" => n11 <= "011010011000110000101101111001011000";
        when "00110010" => n11 <= "011010001010011010101101100100101111";
        when "00110011" => n11 <= "011001111011110100101101010000010010";
        when "00110100" => n11 <= "011001101100111110101100111100000000";
        when "00110101" => n11 <= "011001011101110111101100100111111010";
        when "00110110" => n11 <= "011001001110100010101100010100000000";
        when "00110111" => n11 <= "011000111110111100101100000000010010";
        when "00111000" => n11 <= "011000101111001000101011101100110000";
        when "00111001" => n11 <= "011000011111000100101011011001011011";
        when "00111010" => n11 <= "011000001110110000101011000110010011";
        when "00111011" => n11 <= "010111111110001110101010110011010111";
        when "00111100" => n11 <= "010111101101011101101010100000101001";
        when "00111101" => n11 <= "010111011100011110101010001110001000";
        when "00111110" => n11 <= "010111001011010000101001111011110100";
        when "00111111" => n11 <= "010110111001110100101001101001101110";
        when "01000000" => n11 <= "010110101000001001101001010111110110";
        when "01000001" => n11 <= "010110010110010001101001000110001011";
        when "01000010" => n11 <= "010110000100001011101000110100101111";
        when "01000011" => n11 <= "010101110001110111101000100011100001";
        when "01000100" => n11 <= "010101011111010110101000010010100010";
        when "01000101" => n11 <= "010101001100101000101000000001110001";
        when "01000110" => n11 <= "010100111001101100100111110001001111";
        when "01000111" => n11 <= "010100100110100100100111100000111011";
        when "01001000" => n11 <= "010100010011001111100111010000110111";
        when "01001001" => n11 <= "010011111111101101100111000001000011";
        when "01001010" => n11 <= "010011101011111111100110110001011101";
        when "01001011" => n11 <= "010011011000000101100110100010001000";
        when "01001100" => n11 <= "010011000011111111100110010011000001";
        when "01001101" => n11 <= "010010101111101101100110000100001011";
        when "01001110" => n11 <= "010010011011010000100101110101100101";
        when "01001111" => n11 <= "010010000110100111100101100111001111";
        when "01010000" => n11 <= "010001110001110011100101011001001001";
        when "01010001" => n11 <= "010001011100110100100101001011010100";
        when "01010010" => n11 <= "010001000111101011100100111101101111";
        when "01010011" => n11 <= "010000110010010111100100110000011011";
        when "01010100" => n11 <= "010000011100111000100100100011010111";
        when "01010101" => n11 <= "010000000111001111100100010110100101";
        when "01010110" => n11 <= "001111110001011101100100001010000011";
        when "01010111" => n11 <= "001111011011100000100011111101110011";
        when "01011000" => n11 <= "001111000101011010100011110001110100";
        when "01011001" => n11 <= "001110101111001011100011100110000111";
        when "01011010" => n11 <= "001110011000110011100011011010101011";
        when "01011011" => n11 <= "001110000010010010100011001111100000";
        when "01011100" => n11 <= "001101101011101000100011000100101000";
        when "01011101" => n11 <= "001101010100110110100010111010000001";
        when "01011110" => n11 <= "001100111101111011100010101111101100";
        when "01011111" => n11 <= "001100100110111001100010100101101001";
        when "01100000" => n11 <= "001100001111101111100010011011111001";
        when "01100001" => n11 <= "001011111000011101100010010010011010";
        when "01100010" => n11 <= "001011100001000100100010001001001110";
        when "01100011" => n11 <= "001011001001100011100010000000010101";
        when "01100100" => n11 <= "001010110001111100100001110111101101";
        when "01100101" => n11 <= "001010011010001111100001101111011001";
        when "01100110" => n11 <= "001010000010011010100001100111010111";
        when "01100111" => n11 <= "001001101010100000100001011111101000";
        when "01101000" => n11 <= "001001010010100000100001011000001011";
        when "01101001" => n11 <= "001000111010011010100001010001000010";
        when "01101010" => n11 <= "001000100010001110100001001010001011";
        when "01101011" => n11 <= "001000001001111101100001000011101000";
        when "01101100" => n11 <= "000111110001100111100000111101011000";
        when "01101101" => n11 <= "000111011001001101100000110111011010";
        when "01101110" => n11 <= "000111000000101110100000110001110000";
        when "01101111" => n11 <= "000110101000001010100000101100011001";
        when "01110000" => n11 <= "000110001111100010100000100111010110";
        when "01110001" => n11 <= "000101110110110111100000100010100110";
        when "01110010" => n11 <= "000101011110001000100000011110001001";
        when "01110011" => n11 <= "000101000101010101100000011010000000";
        when "01110100" => n11 <= "000100101100100000100000010110001010";
        when "01110101" => n11 <= "000100010011100111100000010010101000";
        when "01110110" => n11 <= "000011111010101100100000001111011001";
        when "01110111" => n11 <= "000011100001101111100000001100011110";
        when "01111000" => n11 <= "000011001000101111100000001001110111";
        when "01111001" => n11 <= "000010101111101101100000000111100011";
        when "01111010" => n11 <= "000010010110101010100000000101100011";
        when "01111011" => n11 <= "000001111101100101100000000011110110";
        when "01111100" => n11 <= "000001100100011111100000000010011101";
        when "01111101" => n11 <= "000001001011011000100000000001011000";
        when "01111110" => n11 <= "000000110010010000100000000000100111";
        when "01111111" => n11 <= "000000011001001000100000000000001001";
        when "10000000" => n11 <= "000000000000000000100000000000000000";
        when "10000001" => n11 <= "111111100110110111100000000000001001";
        when "10000010" => n11 <= "111111001101101111100000000000100111";
        when "10000011" => n11 <= "111110110100100111100000000001011000";
        when "10000100" => n11 <= "111110011011100000100000000010011101";
        when "10000101" => n11 <= "111110000010011010100000000011110110";
        when "10000110" => n11 <= "111101101001010101100000000101100011";
        when "10000111" => n11 <= "111101010000010010100000000111100011";
        when "10001000" => n11 <= "111100110111010000100000001001110111";
        when "10001001" => n11 <= "111100011110010000100000001100011110";
        when "10001010" => n11 <= "111100000101010011100000001111011001";
        when "10001011" => n11 <= "111011101100011000100000010010101000";
        when "10001100" => n11 <= "111011010011011111100000010110001010";
        when "10001101" => n11 <= "111010111010101010100000011010000000";
        when "10001110" => n11 <= "111010100001110111100000011110001001";
        when "10001111" => n11 <= "111010001001001000100000100010100110";
        when "10010000" => n11 <= "111001110000011101100000100111010110";
        when "10010001" => n11 <= "111001010111110101100000101100011001";
        when "10010010" => n11 <= "111000111111010001100000110001110000";
        when "10010011" => n11 <= "111000100110110010100000110111011010";
        when "10010100" => n11 <= "111000001110011000100000111101011000";
        when "10010101" => n11 <= "110111110110000010100001000011101000";
        when "10010110" => n11 <= "110111011101110001100001001010001011";
        when "10010111" => n11 <= "110111000101100101100001010001000010";
        when "10011000" => n11 <= "110110101101011111100001011000001011";
        when "10011001" => n11 <= "110110010101011111100001011111101000";
        when "10011010" => n11 <= "110101111101100101100001100111010111";
        when "10011011" => n11 <= "110101100101110000100001101111011001";
        when "10011100" => n11 <= "110101001110000011100001110111101101";
        when "10011101" => n11 <= "110100110110011100100010000000010101";
        when "10011110" => n11 <= "110100011110111011100010001001001110";
        when "10011111" => n11 <= "110100000111100010100010010010011010";
        when "10100000" => n11 <= "110011110000010000100010011011111001";
        when "10100001" => n11 <= "110011011001000110100010100101101001";
        when "10100010" => n11 <= "110011000010000100100010101111101100";
        when "10100011" => n11 <= "110010101011001001100010111010000001";
        when "10100100" => n11 <= "110010010100010111100011000100101000";
        when "10100101" => n11 <= "110001111101101101100011001111100000";
        when "10100110" => n11 <= "110001100111001100100011011010101011";
        when "10100111" => n11 <= "110001010000110100100011100110000111";
        when "10101000" => n11 <= "110000111010100101100011110001110100";
        when "10101001" => n11 <= "110000100100011111100011111101110011";
        when "10101010" => n11 <= "110000001110100010100100001010000011";
        when "10101011" => n11 <= "101111111000110000100100010110100101";
        when "10101100" => n11 <= "101111100011000111100100100011010111";
        when "10101101" => n11 <= "101111001101101000100100110000011011";
        when "10101110" => n11 <= "101110111000010100100100111101101111";
        when "10101111" => n11 <= "101110100011001011100101001011010100";
        when "10110000" => n11 <= "101110001110001100100101011001001001";
        when "10110001" => n11 <= "101101111001011000100101100111001111";
        when "10110010" => n11 <= "101101100100101111100101110101100101";
        when "10110011" => n11 <= "101101010000010010100110000100001011";
        when "10110100" => n11 <= "101100111100000000100110010011000001";
        when "10110101" => n11 <= "101100100111111010100110100010001000";
        when "10110110" => n11 <= "101100010100000000100110110001011101";
        when "10110111" => n11 <= "101100000000010010100111000001000011";
        when "10111000" => n11 <= "101011101100110000100111010000110111";
        when "10111001" => n11 <= "101011011001011011100111100000111011";
        when "10111010" => n11 <= "101011000110010011100111110001001111";
        when "10111011" => n11 <= "101010110011010111101000000001110001";
        when "10111100" => n11 <= "101010100000101001101000010010100010";
        when "10111101" => n11 <= "101010001110001000101000100011100001";
        when "10111110" => n11 <= "101001111011110100101000110100101111";
        when "10111111" => n11 <= "101001101001101110101001000110001011";
        when "11000000" => n11 <= "101001010111110110101001010111110110";
        when "11000001" => n11 <= "101001000110001011101001101001101110";
        when "11000010" => n11 <= "101000110100101111101001111011110100";
        when "11000011" => n11 <= "101000100011100001101010001110001000";
        when "11000100" => n11 <= "101000010010100010101010100000101001";
        when "11000101" => n11 <= "101000000001110001101010110011010111";
        when "11000110" => n11 <= "100111110001001111101011000110010011";
        when "11000111" => n11 <= "100111100000111011101011011001011011";
        when "11001000" => n11 <= "100111010000110111101011101100110000";
        when "11001001" => n11 <= "100111000001000011101100000000010010";
        when "11001010" => n11 <= "100110110001011101101100010100000000";
        when "11001011" => n11 <= "100110100010001000101100100111111010";
        when "11001100" => n11 <= "100110010011000001101100111100000000";
        when "11001101" => n11 <= "100110000100001011101101010000010010";
        when "11001110" => n11 <= "100101110101100101101101100100101111";
        when "11001111" => n11 <= "100101100111001111101101111001011000";
        when "11010000" => n11 <= "100101011001001001101110001110001100";
        when "11010001" => n11 <= "100101001011010100101110100011001011";
        when "11010010" => n11 <= "100100111101101111101110111000010100";
        when "11010011" => n11 <= "100100110000011011101111001101101000";
        when "11010100" => n11 <= "100100100011010111101111100011000111";
        when "11010101" => n11 <= "100100010110100101101111111000110000";
        when "11010110" => n11 <= "100100001010000011110000001110100010";
        when "11010111" => n11 <= "100011111101110011110000100100011111";
        when "11011000" => n11 <= "100011110001110100110000111010100101";
        when "11011001" => n11 <= "100011100110000111110001010000110100";
        when "11011010" => n11 <= "100011011010101011110001100111001100";
        when "11011011" => n11 <= "100011001111100000110001111101101101";
        when "11011100" => n11 <= "100011000100101000110010010100010111";
        when "11011101" => n11 <= "100010111010000001110010101011001001";
        when "11011110" => n11 <= "100010101111101100110011000010000100";
        when "11011111" => n11 <= "100010100101101001110011011001000110";
        when "11100000" => n11 <= "100010011011111001110011110000010000";
        when "11100001" => n11 <= "100010010010011010110100000111100010";
        when "11100010" => n11 <= "100010001001001110110100011110111011";
        when "11100011" => n11 <= "100010000000010101110100110110011100";
        when "11100100" => n11 <= "100001110111101101110101001110000011";
        when "11100101" => n11 <= "100001101111011001110101100101110000";
        when "11100110" => n11 <= "100001100111010111110101111101100101";
        when "11100111" => n11 <= "100001011111101000110110010101011111";
        when "11101000" => n11 <= "100001011000001011110110101101011111";
        when "11101001" => n11 <= "100001010001000010110111000101100101";
        when "11101010" => n11 <= "100001001010001011110111011101110001";
        when "11101011" => n11 <= "100001000011101000110111110110000010";
        when "11101100" => n11 <= "100000111101011000111000001110011000";
        when "11101101" => n11 <= "100000110111011010111000100110110010";
        when "11101110" => n11 <= "100000110001110000111000111111010001";
        when "11101111" => n11 <= "100000101100011001111001010111110101";
        when "11110000" => n11 <= "100000100111010110111001110000011101";
        when "11110001" => n11 <= "100000100010100110111010001001001000";
        when "11110010" => n11 <= "100000011110001001111010100001110111";
        when "11110011" => n11 <= "100000011010000000111010111010101010";
        when "11110100" => n11 <= "100000010110001010111011010011011111";
        when "11110101" => n11 <= "100000010010101000111011101100011000";
        when "11110110" => n11 <= "100000001111011001111100000101010011";
        when "11110111" => n11 <= "100000001100011110111100011110010000";
        when "11111000" => n11 <= "100000001001110111111100110111010000";
        when "11111001" => n11 <= "100000000111100011111101010000010010";
        when "11111010" => n11 <= "100000000101100011111101101001010101";
        when "11111011" => n11 <= "100000000011110110111110000010011010";
        when "11111100" => n11 <= "100000000010011101111110011011100000";
        when "11111101" => n11 <= "100000000001011000111110110100100111";
        when "11111110" => n11 <= "100000000000100111111111001101101111";
        when "11111111" => n11 <= "100000000000001001111111100110110111";
        when others => n11 <= "XXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX";
      end case;
    end if;
  end if;
end process;
n12 <= n11(35 downto 35) &
  n11(34 downto 34) &
  n11(33 downto 33) &
  n11(32 downto 32) &
  n11(31 downto 31) &
  n11(30 downto 30) &
  n11(29 downto 29) &
  n11(28 downto 28) &
  n11(27 downto 27) &
  n11(26 downto 26) &
  n11(25 downto 25) &
  n11(24 downto 24) &
  n11(23 downto 23) &
  n11(22 downto 22) &
  n11(21 downto 21) &
  n11(20 downto 20) &
  n11(19 downto 19) &
  n11(18 downto 18);
n13 <= n11(17 downto 17) &
  n11(16 downto 16) &
  n11(15 downto 15) &
  n11(14 downto 14) &
  n11(13 downto 13) &
  n11(12 downto 12) &
  n11(11 downto 11) &
  n11(10 downto 10) &
  n11(9 downto 9) &
  n11(8 downto 8) &
  n11(7 downto 7) &
  n11(6 downto 6) &
  n11(5 downto 5) &
  n11(4 downto 4) &
  n11(3 downto 3) &
  n11(2 downto 2) &
  n11(1 downto 1) &
  n11(0 downto 0);
n14 <= unsigned(signed(n5) * signed(n12));
n15 <= n14(34 downto 34) &
  n14(33 downto 33) &
  n14(32 downto 32) &
  n14(31 downto 31) &
  n14(30 downto 30) &
  n14(29 downto 29) &
  n14(28 downto 28) &
  n14(27 downto 27) &
  n14(26 downto 26) &
  n14(25 downto 25) &
  n14(24 downto 24) &
  n14(23 downto 23) &
  n14(22 downto 22) &
  n14(21 downto 21) &
  n14(20 downto 20) &
  n14(19 downto 19) &
  n14(18 downto 18) &
  n14(17 downto 17);
process (clock_c) begin
  if rising_edge(clock_c) then
    if i5 = "1" then
      n16 <= "000000000000000000";
    elsif i4 = "1" then
      n16 <= n15;
    end if;
  end if;
end process;
n17 <= unsigned(signed(n6) * signed(n13));
n18 <= n17(34 downto 34) &
  n17(33 downto 33) &
  n17(32 downto 32) &
  n17(31 downto 31) &
  n17(30 downto 30) &
  n17(29 downto 29) &
  n17(28 downto 28) &
  n17(27 downto 27) &
  n17(26 downto 26) &
  n17(25 downto 25) &
  n17(24 downto 24) &
  n17(23 downto 23) &
  n17(22 downto 22) &
  n17(21 downto 21) &
  n17(20 downto 20) &
  n17(19 downto 19) &
  n17(18 downto 18) &
  n17(17 downto 17);
process (clock_c) begin
  if rising_edge(clock_c) then
    if i5 = "1" then
      n19 <= "000000000000000000";
    elsif i4 = "1" then
      n19 <= n18;
    end if;
  end if;
end process;
n20 <= n16 - n19;
process (clock_c) begin
  if rising_edge(clock_c) then
    if i5 = "1" then
      n21 <= "000000000000000000";
    elsif i4 = "1" then
      n21 <= n20;
    end if;
  end if;
end process;
n22 <= unsigned(signed(n5) * signed(n13));
n23 <= n22(34 downto 34) &
  n22(33 downto 33) &
  n22(32 downto 32) &
  n22(31 downto 31) &
  n22(30 downto 30) &
  n22(29 downto 29) &
  n22(28 downto 28) &
  n22(27 downto 27) &
  n22(26 downto 26) &
  n22(25 downto 25) &
  n22(24 downto 24) &
  n22(23 downto 23) &
  n22(22 downto 22) &
  n22(21 downto 21) &
  n22(20 downto 20) &
  n22(19 downto 19) &
  n22(18 downto 18) &
  n22(17 downto 17);
process (clock_c) begin
  if rising_edge(clock_c) then
    if i5 = "1" then
      n24 <= "000000000000000000";
    elsif i4 = "1" then
      n24 <= n23;
    end if;
  end if;
end process;
n25 <= unsigned(signed(n6) * signed(n12));
n26 <= n25(34 downto 34) &
  n25(33 downto 33) &
  n25(32 downto 32) &
  n25(31 downto 31) &
  n25(30 downto 30) &
  n25(29 downto 29) &
  n25(28 downto 28) &
  n25(27 downto 27) &
  n25(26 downto 26) &
  n25(25 downto 25) &
  n25(24 downto 24) &
  n25(23 downto 23) &
  n25(22 downto 22) &
  n25(21 downto 21) &
  n25(20 downto 20) &
  n25(19 downto 19) &
  n25(18 downto 18) &
  n25(17 downto 17);
process (clock_c) begin
  if rising_edge(clock_c) then
    if i5 = "1" then
      n27 <= "000000000000000000";
    elsif i4 = "1" then
      n27 <= n26;
    end if;
  end if;
end process;
n28 <= n24 + n27;
process (clock_c) begin
  if rising_edge(clock_c) then
    if i5 = "1" then
      n29 <= "000000000000000000";
    elsif i4 = "1" then
      n29 <= n28;
    end if;
  end if;
end process;
n30 <= n8 + n21;
n31 <= n10 + n29;
n32 <= n30 & n31;
process (clock_c) begin
  if rising_edge(clock_c) then
    if i5 = "1" then
      n33 <= "000000000000000000000000000000000000";
    elsif i4 = "1" then
      n33 <= n32;
    end if;
  end if;
end process;
n34 <= n8 - n21;
n35 <= n10 - n29;
n36 <= n34 & n35;
process (clock_c) begin
  if rising_edge(clock_c) then
    if i5 = "1" then
      n37 <= "000000000000000000000000000000000000";
    elsif i4 = "1" then
      n37 <= n36;
    end if;
  end if;
end process;
o2 <= n37;
o1 <= n33;
end architecture rtl;

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
entity cf_fft_4096_18_19 is
port (
clock_c : in std_logic;
i1 : in  unsigned(0 downto 0);
i2 : in  unsigned(35 downto 0);
i3 : in  unsigned(35 downto 0);
i4 : in  unsigned(0 downto 0);
i5 : in  unsigned(0 downto 0);
o1 : out unsigned(0 downto 0);
o2 : out unsigned(35 downto 0);
o3 : out unsigned(35 downto 0));
end entity cf_fft_4096_18_19;
architecture rtl of cf_fft_4096_18_19 is
signal n1 : unsigned(7 downto 0);
signal n2 : unsigned(71 downto 0);
signal n3 : unsigned(0 downto 0) := "0";
signal n4 : unsigned(0 downto 0) := "0";
signal n5 : unsigned(0 downto 0) := "0";
signal n6 : unsigned(0 downto 0) := "0";
signal n7 : unsigned(9 downto 0);
signal n8 : unsigned(9 downto 0) := "0000000000";
signal n9 : unsigned(9 downto 0) := "0000000000";
signal n10 : unsigned(9 downto 0) := "0000000000";
signal n11 : unsigned(9 downto 0) := "0000000000";
signal n12 : unsigned(0 downto 0);
signal n13 : unsigned(0 downto 0) := "0";
signal n14 : unsigned(0 downto 0) := "0";
signal n15 : unsigned(0 downto 0) := "0";
signal n16 : unsigned(0 downto 0) := "0";
signal n17 : unsigned(0 downto 0);
signal n18 : unsigned(1 downto 0);
signal n19 : unsigned(35 downto 0);
signal n20 : unsigned(35 downto 0);
signal n21 : unsigned(35 downto 0);
signal n22 : unsigned(35 downto 0);
signal n23 : unsigned(35 downto 0);
signal n24 : unsigned(35 downto 0);
signal s25_1 : unsigned(35 downto 0);
signal s25_2 : unsigned(35 downto 0);
signal s26_1 : unsigned(0 downto 0);
signal s27_1 : unsigned(71 downto 0);
signal s28_1 : unsigned(0 downto 0);
signal s28_2 : unsigned(0 downto 0);
signal s28_3 : unsigned(71 downto 0);
signal s29_1 : unsigned(10 downto 0);
signal s29_2 : unsigned(0 downto 0);
component cf_fft_4096_18_20 is
port (
clock_c : in std_logic;
i1 : in  unsigned(35 downto 0);
i2 : in  unsigned(35 downto 0);
i3 : in  unsigned(7 downto 0);
i4 : in  unsigned(0 downto 0);
i5 : in  unsigned(0 downto 0);
o1 : out unsigned(35 downto 0);
o2 : out unsigned(35 downto 0));
end component cf_fft_4096_18_20;
component cf_fft_4096_18_37 is
port (
clock_c : in std_logic;
i1 : in  unsigned(1 downto 0);
i2 : in  unsigned(0 downto 0);
i3 : in  unsigned(0 downto 0);
o1 : out unsigned(0 downto 0));
end component cf_fft_4096_18_37;
component cf_fft_4096_18_33 is
port (
clock_c : in std_logic;
i1 : in  unsigned(71 downto 0);
i2 : in  unsigned(0 downto 0);
i3 : in  unsigned(9 downto 0);
i4 : in  unsigned(0 downto 0);
i5 : in  unsigned(0 downto 0);
i6 : in  unsigned(0 downto 0);
o1 : out unsigned(71 downto 0));
end component cf_fft_4096_18_33;
component cf_fft_4096_18_32 is
port (
clock_c : in std_logic;
i1 : in  unsigned(71 downto 0);
i2 : in  unsigned(0 downto 0);
i3 : in  unsigned(9 downto 0);
i4 : in  unsigned(0 downto 0);
i5 : in  unsigned(0 downto 0);
i6 : in  unsigned(0 downto 0);
o1 : out unsigned(0 downto 0);
o2 : out unsigned(0 downto 0);
o3 : out unsigned(71 downto 0));
end component cf_fft_4096_18_32;
component cf_fft_4096_18_28 is
port (
clock_c : in std_logic;
i1 : in  unsigned(0 downto 0);
i2 : in  unsigned(0 downto 0);
i3 : in  unsigned(0 downto 0);
o1 : out unsigned(10 downto 0);
o2 : out unsigned(0 downto 0));
end component cf_fft_4096_18_28;
begin
n1 <= s29_1(10 downto 10) &
  s29_1(9 downto 9) &
  s29_1(8 downto 8) &
  s29_1(7 downto 7) &
  s29_1(6 downto 6) &
  s29_1(5 downto 5) &
  s29_1(4 downto 4) &
  s29_1(3 downto 3);
n2 <= s25_1 & s25_2;
process (clock_c) begin
  if rising_edge(clock_c) then
    if i5 = "1" then
      n3 <= "0";
    elsif i4 = "1" then
      n3 <= s29_2;
    end if;
  end if;
end process;
process (clock_c) begin
  if rising_edge(clock_c) then
    if i5 = "1" then
      n4 <= "0";
    elsif i4 = "1" then
      n4 <= n3;
    end if;
  end if;
end process;
process (clock_c) begin
  if rising_edge(clock_c) then
    if i5 = "1" then
      n5 <= "0";
    elsif i4 = "1" then
      n5 <= n4;
    end if;
  end if;
end process;
process (clock_c) begin
  if rising_edge(clock_c) then
    if i5 = "1" then
      n6 <= "0";
    elsif i4 = "1" then
      n6 <= n5;
    end if;
  end if;
end process;
n7 <= s29_1(10 downto 10) &
  s29_1(9 downto 9) &
  s29_1(8 downto 8) &
  s29_1(7 downto 7) &
  s29_1(6 downto 6) &
  s29_1(5 downto 5) &
  s29_1(4 downto 4) &
  s29_1(3 downto 3) &
  s29_1(2 downto 2) &
  s29_1(1 downto 1);
process (clock_c) begin
  if rising_edge(clock_c) then
    if i5 = "1" then
      n8 <= "0000000000";
    elsif i4 = "1" then
      n8 <= n7;
    end if;
  end if;
end process;
process (clock_c) begin
  if rising_edge(clock_c) then
    if i5 = "1" then
      n9 <= "0000000000";
    elsif i4 = "1" then
      n9 <= n8;
    end if;
  end if;
end process;
process (clock_c) begin
  if rising_edge(clock_c) then
    if i5 = "1" then
      n10 <= "0000000000";
    elsif i4 = "1" then
      n10 <= n9;
    end if;
  end if;
end process;
process (clock_c) begin
  if rising_edge(clock_c) then
    if i5 = "1" then
      n11 <= "0000000000";
    elsif i4 = "1" then
      n11 <= n10;
    end if;
  end if;
end process;
n12 <= s29_1(0 downto 0);
process (clock_c) begin
  if rising_edge(clock_c) then
    if i5 = "1" then
      n13 <= "0";
    elsif i4 = "1" then
      n13 <= n12;
    end if;
  end if;
end process;
process (clock_c) begin
  if rising_edge(clock_c) then
    if i5 = "1" then
      n14 <= "0";
    elsif i4 = "1" then
      n14 <= n13;
    end if;
  end if;
end process;
process (clock_c) begin
  if rising_edge(clock_c) then
    if i5 = "1" then
      n15 <= "0";
    elsif i4 = "1" then
      n15 <= n14;
    end if;
  end if;
end process;
process (clock_c) begin
  if rising_edge(clock_c) then
    if i5 = "1" then
      n16 <= "0";
    elsif i4 = "1" then
      n16 <= n15;
    end if;
  end if;
end process;
n17 <= not n16;
n18 <= s28_2 & s28_1;
n19 <= s28_3(71 downto 71) &
  s28_3(70 downto 70) &
  s28_3(69 downto 69) &
  s28_3(68 downto 68) &
  s28_3(67 downto 67) &
  s28_3(66 downto 66) &
  s28_3(65 downto 65) &
  s28_3(64 downto 64) &
  s28_3(63 downto 63) &
  s28_3(62 downto 62) &
  s28_3(61 downto 61) &
  s28_3(60 downto 60) &
  s28_3(59 downto 59) &
  s28_3(58 downto 58) &
  s28_3(57 downto 57) &
  s28_3(56 downto 56) &
  s28_3(55 downto 55) &
  s28_3(54 downto 54) &
  s28_3(53 downto 53) &
  s28_3(52 downto 52) &
  s28_3(51 downto 51) &
  s28_3(50 downto 50) &
  s28_3(49 downto 49) &
  s28_3(48 downto 48) &
  s28_3(47 downto 47) &
  s28_3(46 downto 46) &
  s28_3(45 downto 45) &
  s28_3(44 downto 44) &
  s28_3(43 downto 43) &
  s28_3(42 downto 42) &
  s28_3(41 downto 41) &
  s28_3(40 downto 40) &
  s28_3(39 downto 39) &
  s28_3(38 downto 38) &
  s28_3(37 downto 37) &
  s28_3(36 downto 36);
n20 <= s28_3(35 downto 35) &
  s28_3(34 downto 34) &
  s28_3(33 downto 33) &
  s28_3(32 downto 32) &
  s28_3(31 downto 31) &
  s28_3(30 downto 30) &
  s28_3(29 downto 29) &
  s28_3(28 downto 28) &
  s28_3(27 downto 27) &
  s28_3(26 downto 26) &
  s28_3(25 downto 25) &
  s28_3(24 downto 24) &
  s28_3(23 downto 23) &
  s28_3(22 downto 22) &
  s28_3(21 downto 21) &
  s28_3(20 downto 20) &
  s28_3(19 downto 19) &
  s28_3(18 downto 18) &
  s28_3(17 downto 17) &
  s28_3(16 downto 16) &
  s28_3(15 downto 15) &
  s28_3(14 downto 14) &
  s28_3(13 downto 13) &
  s28_3(12 downto 12) &
  s28_3(11 downto 11) &
  s28_3(10 downto 10) &
  s28_3(9 downto 9) &
  s28_3(8 downto 8) &
  s28_3(7 downto 7) &
  s28_3(6 downto 6) &
  s28_3(5 downto 5) &
  s28_3(4 downto 4) &
  s28_3(3 downto 3) &
  s28_3(2 downto 2) &
  s28_3(1 downto 1) &
  s28_3(0 downto 0);
n21 <= s27_1(71 downto 71) &
  s27_1(70 downto 70) &
  s27_1(69 downto 69) &
  s27_1(68 downto 68) &
  s27_1(67 downto 67) &
  s27_1(66 downto 66) &
  s27_1(65 downto 65) &
  s27_1(64 downto 64) &
  s27_1(63 downto 63) &
  s27_1(62 downto 62) &
  s27_1(61 downto 61) &
  s27_1(60 downto 60) &
  s27_1(59 downto 59) &
  s27_1(58 downto 58) &
  s27_1(57 downto 57) &
  s27_1(56 downto 56) &
  s27_1(55 downto 55) &
  s27_1(54 downto 54) &
  s27_1(53 downto 53) &
  s27_1(52 downto 52) &
  s27_1(51 downto 51) &
  s27_1(50 downto 50) &
  s27_1(49 downto 49) &
  s27_1(48 downto 48) &
  s27_1(47 downto 47) &
  s27_1(46 downto 46) &
  s27_1(45 downto 45) &
  s27_1(44 downto 44) &
  s27_1(43 downto 43) &
  s27_1(42 downto 42) &
  s27_1(41 downto 41) &
  s27_1(40 downto 40) &
  s27_1(39 downto 39) &
  s27_1(38 downto 38) &
  s27_1(37 downto 37) &
  s27_1(36 downto 36);
n22 <= s27_1(35 downto 35) &
  s27_1(34 downto 34) &
  s27_1(33 downto 33) &
  s27_1(32 downto 32) &
  s27_1(31 downto 31) &
  s27_1(30 downto 30) &
  s27_1(29 downto 29) &
  s27_1(28 downto 28) &
  s27_1(27 downto 27) &
  s27_1(26 downto 26) &
  s27_1(25 downto 25) &
  s27_1(24 downto 24) &
  s27_1(23 downto 23) &
  s27_1(22 downto 22) &
  s27_1(21 downto 21) &
  s27_1(20 downto 20) &
  s27_1(19 downto 19) &
  s27_1(18 downto 18) &
  s27_1(17 downto 17) &
  s27_1(16 downto 16) &
  s27_1(15 downto 15) &
  s27_1(14 downto 14) &
  s27_1(13 downto 13) &
  s27_1(12 downto 12) &
  s27_1(11 downto 11) &
  s27_1(10 downto 10) &
  s27_1(9 downto 9) &
  s27_1(8 downto 8) &
  s27_1(7 downto 7) &
  s27_1(6 downto 6) &
  s27_1(5 downto 5) &
  s27_1(4 downto 4) &
  s27_1(3 downto 3) &
  s27_1(2 downto 2) &
  s27_1(1 downto 1) &
  s27_1(0 downto 0);
n23 <= n20 when s26_1 = "1" else n19;
n24 <= n22 when s26_1 = "1" else n21;
s25 : cf_fft_4096_18_20 port map (clock_c, i2, i3, n1, i4, i5, s25_1, s25_2);
s26 : cf_fft_4096_18_37 port map (clock_c, n18, i4, i5, s26_1);
s27 : cf_fft_4096_18_33 port map (clock_c, n2, n6, n11, n16, i4, i5, s27_1);
s28 : cf_fft_4096_18_32 port map (clock_c, n2, n6, n11, n17, i4, i5, s28_1, s28_2, s28_3);
s29 : cf_fft_4096_18_28 port map (clock_c, i1, i4, i5, s29_1, s29_2);
o3 <= n24;
o2 <= n23;
o1 <= s28_1;
end architecture rtl;

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
entity cf_fft_4096_18_18 is
port (
clock_c : in std_logic;
i1 : in  unsigned(35 downto 0);
i2 : in  unsigned(35 downto 0);
i3 : in  unsigned(6 downto 0);
i4 : in  unsigned(0 downto 0);
i5 : in  unsigned(0 downto 0);
o1 : out unsigned(35 downto 0);
o2 : out unsigned(35 downto 0));
end entity cf_fft_4096_18_18;
architecture rtl of cf_fft_4096_18_18 is
signal n1 : unsigned(35 downto 0) := "000000000000000000000000000000000000";
signal n2 : unsigned(17 downto 0);
signal n3 : unsigned(17 downto 0);
signal n4 : unsigned(35 downto 0) := "000000000000000000000000000000000000";
signal n5 : unsigned(17 downto 0);
signal n6 : unsigned(17 downto 0);
signal n7 : unsigned(17 downto 0) := "000000000000000000";
signal n8 : unsigned(17 downto 0) := "000000000000000000";
signal n9 : unsigned(17 downto 0) := "000000000000000000";
signal n10 : unsigned(17 downto 0) := "000000000000000000";
signal n11 : unsigned(35 downto 0) := "000000000000000000000000000000000000";
signal n12 : unsigned(17 downto 0);
signal n13 : unsigned(17 downto 0);
signal n14 : unsigned(35 downto 0);
signal n15 : unsigned(17 downto 0);
signal n16 : unsigned(17 downto 0) := "000000000000000000";
signal n17 : unsigned(35 downto 0);
signal n18 : unsigned(17 downto 0);
signal n19 : unsigned(17 downto 0) := "000000000000000000";
signal n20 : unsigned(17 downto 0);
signal n21 : unsigned(17 downto 0) := "000000000000000000";
signal n22 : unsigned(35 downto 0);
signal n23 : unsigned(17 downto 0);
signal n24 : unsigned(17 downto 0) := "000000000000000000";
signal n25 : unsigned(35 downto 0);
signal n26 : unsigned(17 downto 0);
signal n27 : unsigned(17 downto 0) := "000000000000000000";
signal n28 : unsigned(17 downto 0);
signal n29 : unsigned(17 downto 0) := "000000000000000000";
signal n30 : unsigned(17 downto 0);
signal n31 : unsigned(17 downto 0);
signal n32 : unsigned(35 downto 0);
signal n33 : unsigned(35 downto 0) := "000000000000000000000000000000000000";
signal n34 : unsigned(17 downto 0);
signal n35 : unsigned(17 downto 0);
signal n36 : unsigned(35 downto 0);
signal n37 : unsigned(35 downto 0) := "000000000000000000000000000000000000";
begin
process (clock_c) begin
  if rising_edge(clock_c) then
    if i5 = "1" then
      n1 <= "000000000000000000000000000000000000";
    elsif i4 = "1" then
      n1 <= i1;
    end if;
  end if;
end process;
n2 <= n1(35 downto 35) &
  n1(34 downto 34) &
  n1(33 downto 33) &
  n1(32 downto 32) &
  n1(31 downto 31) &
  n1(30 downto 30) &
  n1(29 downto 29) &
  n1(28 downto 28) &
  n1(27 downto 27) &
  n1(26 downto 26) &
  n1(25 downto 25) &
  n1(24 downto 24) &
  n1(23 downto 23) &
  n1(22 downto 22) &
  n1(21 downto 21) &
  n1(20 downto 20) &
  n1(19 downto 19) &
  n1(18 downto 18);
n3 <= n1(17 downto 17) &
  n1(16 downto 16) &
  n1(15 downto 15) &
  n1(14 downto 14) &
  n1(13 downto 13) &
  n1(12 downto 12) &
  n1(11 downto 11) &
  n1(10 downto 10) &
  n1(9 downto 9) &
  n1(8 downto 8) &
  n1(7 downto 7) &
  n1(6 downto 6) &
  n1(5 downto 5) &
  n1(4 downto 4) &
  n1(3 downto 3) &
  n1(2 downto 2) &
  n1(1 downto 1) &
  n1(0 downto 0);
process (clock_c) begin
  if rising_edge(clock_c) then
    if i5 = "1" then
      n4 <= "000000000000000000000000000000000000";
    elsif i4 = "1" then
      n4 <= i2;
    end if;
  end if;
end process;
n5 <= n4(35 downto 35) &
  n4(34 downto 34) &
  n4(33 downto 33) &
  n4(32 downto 32) &
  n4(31 downto 31) &
  n4(30 downto 30) &
  n4(29 downto 29) &
  n4(28 downto 28) &
  n4(27 downto 27) &
  n4(26 downto 26) &
  n4(25 downto 25) &
  n4(24 downto 24) &
  n4(23 downto 23) &
  n4(22 downto 22) &
  n4(21 downto 21) &
  n4(20 downto 20) &
  n4(19 downto 19) &
  n4(18 downto 18);
n6 <= n4(17 downto 17) &
  n4(16 downto 16) &
  n4(15 downto 15) &
  n4(14 downto 14) &
  n4(13 downto 13) &
  n4(12 downto 12) &
  n4(11 downto 11) &
  n4(10 downto 10) &
  n4(9 downto 9) &
  n4(8 downto 8) &
  n4(7 downto 7) &
  n4(6 downto 6) &
  n4(5 downto 5) &
  n4(4 downto 4) &
  n4(3 downto 3) &
  n4(2 downto 2) &
  n4(1 downto 1) &
  n4(0 downto 0);
process (clock_c) begin
  if rising_edge(clock_c) then
    if i5 = "1" then
      n7 <= "000000000000000000";
    elsif i4 = "1" then
      n7 <= n2;
    end if;
  end if;
end process;
process (clock_c) begin
  if rising_edge(clock_c) then
    if i5 = "1" then
      n8 <= "000000000000000000";
    elsif i4 = "1" then
      n8 <= n7;
    end if;
  end if;
end process;
process (clock_c) begin
  if rising_edge(clock_c) then
    if i5 = "1" then
      n9 <= "000000000000000000";
    elsif i4 = "1" then
      n9 <= n3;
    end if;
  end if;
end process;
process (clock_c) begin
  if rising_edge(clock_c) then
    if i5 = "1" then
      n10 <= "000000000000000000";
    elsif i4 = "1" then
      n10 <= n9;
    end if;
  end if;
end process;
process (clock_c) begin
  if rising_edge(clock_c) then 
    if i4 = "1" then
      case i3 is
        when "0000000" => n11 <= "011111111111111111000000000000000000";
        when "0000001" => n11 <= "011111111111011000111111001101101111";
        when "0000010" => n11 <= "011111111101100010111110011011100000";
        when "0000011" => n11 <= "011111111010011100111101101001010101";
        when "0000100" => n11 <= "011111110110001000111100110111010000";
        when "0000101" => n11 <= "011111110000100110111100000101010011";
        when "0000110" => n11 <= "011111101001110101111011010011011111";
        when "0000111" => n11 <= "011111100001110110111010100001110111";
        when "0001000" => n11 <= "011111011000101001111001110000011101";
        when "0001001" => n11 <= "011111001110001111111000111111010001";
        when "0001010" => n11 <= "011111000010100111111000001110011000";
        when "0001011" => n11 <= "011110110101110100110111011101110001";
        when "0001100" => n11 <= "011110100111110100110110101101011111";
        when "0001101" => n11 <= "011110011000101000110101111101100101";
        when "0001110" => n11 <= "011110001000010010110101001110000011";
        when "0001111" => n11 <= "011101110110110001110100011110111011";
        when "0010000" => n11 <= "011101100100000110110011110000010000";
        when "0010001" => n11 <= "011101010000010011110011000010000100";
        when "0010010" => n11 <= "011100111011010111110010010100010111";
        when "0010011" => n11 <= "011100100101010100110001100111001100";
        when "0010100" => n11 <= "011100001110001011110000111010100101";
        when "0010101" => n11 <= "011011110101111100110000001110100010";
        when "0010110" => n11 <= "011011011100101000101111100011000111";
        when "0010111" => n11 <= "011011000010010000101110111000010100";
        when "0011000" => n11 <= "011010100110110110101110001110001100";
        when "0011001" => n11 <= "011010001010011010101101100100101111";
        when "0011010" => n11 <= "011001101100111110101100111100000000";
        when "0011011" => n11 <= "011001001110100010101100010100000000";
        when "0011100" => n11 <= "011000101111001000101011101100110000";
        when "0011101" => n11 <= "011000001110110000101011000110010011";
        when "0011110" => n11 <= "010111101101011101101010100000101001";
        when "0011111" => n11 <= "010111001011010000101001111011110100";
        when "0100000" => n11 <= "010110101000001001101001010111110110";
        when "0100001" => n11 <= "010110000100001011101000110100101111";
        when "0100010" => n11 <= "010101011111010110101000010010100010";
        when "0100011" => n11 <= "010100111001101100100111110001001111";
        when "0100100" => n11 <= "010100010011001111100111010000110111";
        when "0100101" => n11 <= "010011101011111111100110110001011101";
        when "0100110" => n11 <= "010011000011111111100110010011000001";
        when "0100111" => n11 <= "010010011011010000100101110101100101";
        when "0101000" => n11 <= "010001110001110011100101011001001001";
        when "0101001" => n11 <= "010001000111101011100100111101101111";
        when "0101010" => n11 <= "010000011100111000100100100011010111";
        when "0101011" => n11 <= "001111110001011101100100001010000011";
        when "0101100" => n11 <= "001111000101011010100011110001110100";
        when "0101101" => n11 <= "001110011000110011100011011010101011";
        when "0101110" => n11 <= "001101101011101000100011000100101000";
        when "0101111" => n11 <= "001100111101111011100010101111101100";
        when "0110000" => n11 <= "001100001111101111100010011011111001";
        when "0110001" => n11 <= "001011100001000100100010001001001110";
        when "0110010" => n11 <= "001010110001111100100001110111101101";
        when "0110011" => n11 <= "001010000010011010100001100111010111";
        when "0110100" => n11 <= "001001010010100000100001011000001011";
        when "0110101" => n11 <= "001000100010001110100001001010001011";
        when "0110110" => n11 <= "000111110001100111100000111101011000";
        when "0110111" => n11 <= "000111000000101110100000110001110000";
        when "0111000" => n11 <= "000110001111100010100000100111010110";
        when "0111001" => n11 <= "000101011110001000100000011110001001";
        when "0111010" => n11 <= "000100101100100000100000010110001010";
        when "0111011" => n11 <= "000011111010101100100000001111011001";
        when "0111100" => n11 <= "000011001000101111100000001001110111";
        when "0111101" => n11 <= "000010010110101010100000000101100011";
        when "0111110" => n11 <= "000001100100011111100000000010011101";
        when "0111111" => n11 <= "000000110010010000100000000000100111";
        when "1000000" => n11 <= "000000000000000000100000000000000000";
        when "1000001" => n11 <= "111111001101101111100000000000100111";
        when "1000010" => n11 <= "111110011011100000100000000010011101";
        when "1000011" => n11 <= "111101101001010101100000000101100011";
        when "1000100" => n11 <= "111100110111010000100000001001110111";
        when "1000101" => n11 <= "111100000101010011100000001111011001";
        when "1000110" => n11 <= "111011010011011111100000010110001010";
        when "1000111" => n11 <= "111010100001110111100000011110001001";
        when "1001000" => n11 <= "111001110000011101100000100111010110";
        when "1001001" => n11 <= "111000111111010001100000110001110000";
        when "1001010" => n11 <= "111000001110011000100000111101011000";
        when "1001011" => n11 <= "110111011101110001100001001010001011";
        when "1001100" => n11 <= "110110101101011111100001011000001011";
        when "1001101" => n11 <= "110101111101100101100001100111010111";
        when "1001110" => n11 <= "110101001110000011100001110111101101";
        when "1001111" => n11 <= "110100011110111011100010001001001110";
        when "1010000" => n11 <= "110011110000010000100010011011111001";
        when "1010001" => n11 <= "110011000010000100100010101111101100";
        when "1010010" => n11 <= "110010010100010111100011000100101000";
        when "1010011" => n11 <= "110001100111001100100011011010101011";
        when "1010100" => n11 <= "110000111010100101100011110001110100";
        when "1010101" => n11 <= "110000001110100010100100001010000011";
        when "1010110" => n11 <= "101111100011000111100100100011010111";
        when "1010111" => n11 <= "101110111000010100100100111101101111";
        when "1011000" => n11 <= "101110001110001100100101011001001001";
        when "1011001" => n11 <= "101101100100101111100101110101100101";
        when "1011010" => n11 <= "101100111100000000100110010011000001";
        when "1011011" => n11 <= "101100010100000000100110110001011101";
        when "1011100" => n11 <= "101011101100110000100111010000110111";
        when "1011101" => n11 <= "101011000110010011100111110001001111";
        when "1011110" => n11 <= "101010100000101001101000010010100010";
        when "1011111" => n11 <= "101001111011110100101000110100101111";
        when "1100000" => n11 <= "101001010111110110101001010111110110";
        when "1100001" => n11 <= "101000110100101111101001111011110100";
        when "1100010" => n11 <= "101000010010100010101010100000101001";
        when "1100011" => n11 <= "100111110001001111101011000110010011";
        when "1100100" => n11 <= "100111010000110111101011101100110000";
        when "1100101" => n11 <= "100110110001011101101100010100000000";
        when "1100110" => n11 <= "100110010011000001101100111100000000";
        when "1100111" => n11 <= "100101110101100101101101100100101111";
        when "1101000" => n11 <= "100101011001001001101110001110001100";
        when "1101001" => n11 <= "100100111101101111101110111000010100";
        when "1101010" => n11 <= "100100100011010111101111100011000111";
        when "1101011" => n11 <= "100100001010000011110000001110100010";
        when "1101100" => n11 <= "100011110001110100110000111010100101";
        when "1101101" => n11 <= "100011011010101011110001100111001100";
        when "1101110" => n11 <= "100011000100101000110010010100010111";
        when "1101111" => n11 <= "100010101111101100110011000010000100";
        when "1110000" => n11 <= "100010011011111001110011110000010000";
        when "1110001" => n11 <= "100010001001001110110100011110111011";
        when "1110010" => n11 <= "100001110111101101110101001110000011";
        when "1110011" => n11 <= "100001100111010111110101111101100101";
        when "1110100" => n11 <= "100001011000001011110110101101011111";
        when "1110101" => n11 <= "100001001010001011110111011101110001";
        when "1110110" => n11 <= "100000111101011000111000001110011000";
        when "1110111" => n11 <= "100000110001110000111000111111010001";
        when "1111000" => n11 <= "100000100111010110111001110000011101";
        when "1111001" => n11 <= "100000011110001001111010100001110111";
        when "1111010" => n11 <= "100000010110001010111011010011011111";
        when "1111011" => n11 <= "100000001111011001111100000101010011";
        when "1111100" => n11 <= "100000001001110111111100110111010000";
        when "1111101" => n11 <= "100000000101100011111101101001010101";
        when "1111110" => n11 <= "100000000010011101111110011011100000";
        when "1111111" => n11 <= "100000000000100111111111001101101111";
        when others => n11 <= "XXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX";
      end case;
    end if;
  end if;
end process;
n12 <= n11(35 downto 35) &
  n11(34 downto 34) &
  n11(33 downto 33) &
  n11(32 downto 32) &
  n11(31 downto 31) &
  n11(30 downto 30) &
  n11(29 downto 29) &
  n11(28 downto 28) &
  n11(27 downto 27) &
  n11(26 downto 26) &
  n11(25 downto 25) &
  n11(24 downto 24) &
  n11(23 downto 23) &
  n11(22 downto 22) &
  n11(21 downto 21) &
  n11(20 downto 20) &
  n11(19 downto 19) &
  n11(18 downto 18);
n13 <= n11(17 downto 17) &
  n11(16 downto 16) &
  n11(15 downto 15) &
  n11(14 downto 14) &
  n11(13 downto 13) &
  n11(12 downto 12) &
  n11(11 downto 11) &
  n11(10 downto 10) &
  n11(9 downto 9) &
  n11(8 downto 8) &
  n11(7 downto 7) &
  n11(6 downto 6) &
  n11(5 downto 5) &
  n11(4 downto 4) &
  n11(3 downto 3) &
  n11(2 downto 2) &
  n11(1 downto 1) &
  n11(0 downto 0);
n14 <= unsigned(signed(n5) * signed(n12));
n15 <= n14(34 downto 34) &
  n14(33 downto 33) &
  n14(32 downto 32) &
  n14(31 downto 31) &
  n14(30 downto 30) &
  n14(29 downto 29) &
  n14(28 downto 28) &
  n14(27 downto 27) &
  n14(26 downto 26) &
  n14(25 downto 25) &
  n14(24 downto 24) &
  n14(23 downto 23) &
  n14(22 downto 22) &
  n14(21 downto 21) &
  n14(20 downto 20) &
  n14(19 downto 19) &
  n14(18 downto 18) &
  n14(17 downto 17);
process (clock_c) begin
  if rising_edge(clock_c) then
    if i5 = "1" then
      n16 <= "000000000000000000";
    elsif i4 = "1" then
      n16 <= n15;
    end if;
  end if;
end process;
n17 <= unsigned(signed(n6) * signed(n13));
n18 <= n17(34 downto 34) &
  n17(33 downto 33) &
  n17(32 downto 32) &
  n17(31 downto 31) &
  n17(30 downto 30) &
  n17(29 downto 29) &
  n17(28 downto 28) &
  n17(27 downto 27) &
  n17(26 downto 26) &
  n17(25 downto 25) &
  n17(24 downto 24) &
  n17(23 downto 23) &
  n17(22 downto 22) &
  n17(21 downto 21) &
  n17(20 downto 20) &
  n17(19 downto 19) &
  n17(18 downto 18) &
  n17(17 downto 17);
process (clock_c) begin
  if rising_edge(clock_c) then
    if i5 = "1" then
      n19 <= "000000000000000000";
    elsif i4 = "1" then
      n19 <= n18;
    end if;
  end if;
end process;
n20 <= n16 - n19;
process (clock_c) begin
  if rising_edge(clock_c) then
    if i5 = "1" then
      n21 <= "000000000000000000";
    elsif i4 = "1" then
      n21 <= n20;
    end if;
  end if;
end process;
n22 <= unsigned(signed(n5) * signed(n13));
n23 <= n22(34 downto 34) &
  n22(33 downto 33) &
  n22(32 downto 32) &
  n22(31 downto 31) &
  n22(30 downto 30) &
  n22(29 downto 29) &
  n22(28 downto 28) &
  n22(27 downto 27) &
  n22(26 downto 26) &
  n22(25 downto 25) &
  n22(24 downto 24) &
  n22(23 downto 23) &
  n22(22 downto 22) &
  n22(21 downto 21) &
  n22(20 downto 20) &
  n22(19 downto 19) &
  n22(18 downto 18) &
  n22(17 downto 17);
process (clock_c) begin
  if rising_edge(clock_c) then
    if i5 = "1" then
      n24 <= "000000000000000000";
    elsif i4 = "1" then
      n24 <= n23;
    end if;
  end if;
end process;
n25 <= unsigned(signed(n6) * signed(n12));
n26 <= n25(34 downto 34) &
  n25(33 downto 33) &
  n25(32 downto 32) &
  n25(31 downto 31) &
  n25(30 downto 30) &
  n25(29 downto 29) &
  n25(28 downto 28) &
  n25(27 downto 27) &
  n25(26 downto 26) &
  n25(25 downto 25) &
  n25(24 downto 24) &
  n25(23 downto 23) &
  n25(22 downto 22) &
  n25(21 downto 21) &
  n25(20 downto 20) &
  n25(19 downto 19) &
  n25(18 downto 18) &
  n25(17 downto 17);
process (clock_c) begin
  if rising_edge(clock_c) then
    if i5 = "1" then
      n27 <= "000000000000000000";
    elsif i4 = "1" then
      n27 <= n26;
    end if;
  end if;
end process;
n28 <= n24 + n27;
process (clock_c) begin
  if rising_edge(clock_c) then
    if i5 = "1" then
      n29 <= "000000000000000000";
    elsif i4 = "1" then
      n29 <= n28;
    end if;
  end if;
end process;
n30 <= n8 + n21;
n31 <= n10 + n29;
n32 <= n30 & n31;
process (clock_c) begin
  if rising_edge(clock_c) then
    if i5 = "1" then
      n33 <= "000000000000000000000000000000000000";
    elsif i4 = "1" then
      n33 <= n32;
    end if;
  end if;
end process;
n34 <= n8 - n21;
n35 <= n10 - n29;
n36 <= n34 & n35;
process (clock_c) begin
  if rising_edge(clock_c) then
    if i5 = "1" then
      n37 <= "000000000000000000000000000000000000";
    elsif i4 = "1" then
      n37 <= n36;
    end if;
  end if;
end process;
o2 <= n37;
o1 <= n33;
end architecture rtl;

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
entity cf_fft_4096_18_17 is
port (
clock_c : in std_logic;
i1 : in  unsigned(0 downto 0);
i2 : in  unsigned(35 downto 0);
i3 : in  unsigned(35 downto 0);
i4 : in  unsigned(0 downto 0);
i5 : in  unsigned(0 downto 0);
o1 : out unsigned(0 downto 0);
o2 : out unsigned(35 downto 0);
o3 : out unsigned(35 downto 0));
end entity cf_fft_4096_18_17;
architecture rtl of cf_fft_4096_18_17 is
signal n1 : unsigned(6 downto 0);
signal n2 : unsigned(71 downto 0);
signal n3 : unsigned(0 downto 0) := "0";
signal n4 : unsigned(0 downto 0) := "0";
signal n5 : unsigned(0 downto 0) := "0";
signal n6 : unsigned(0 downto 0) := "0";
signal n7 : unsigned(9 downto 0);
signal n8 : unsigned(9 downto 0) := "0000000000";
signal n9 : unsigned(9 downto 0) := "0000000000";
signal n10 : unsigned(9 downto 0) := "0000000000";
signal n11 : unsigned(9 downto 0) := "0000000000";
signal n12 : unsigned(0 downto 0);
signal n13 : unsigned(0 downto 0) := "0";
signal n14 : unsigned(0 downto 0) := "0";
signal n15 : unsigned(0 downto 0) := "0";
signal n16 : unsigned(0 downto 0) := "0";
signal n17 : unsigned(0 downto 0);
signal n18 : unsigned(1 downto 0);
signal n19 : unsigned(35 downto 0);
signal n20 : unsigned(35 downto 0);
signal n21 : unsigned(35 downto 0);
signal n22 : unsigned(35 downto 0);
signal n23 : unsigned(35 downto 0);
signal n24 : unsigned(35 downto 0);
signal s25_1 : unsigned(35 downto 0);
signal s25_2 : unsigned(35 downto 0);
signal s26_1 : unsigned(0 downto 0);
signal s27_1 : unsigned(10 downto 0);
signal s27_2 : unsigned(0 downto 0);
signal s28_1 : unsigned(71 downto 0);
signal s29_1 : unsigned(0 downto 0);
signal s29_2 : unsigned(0 downto 0);
signal s29_3 : unsigned(71 downto 0);
component cf_fft_4096_18_18 is
port (
clock_c : in std_logic;
i1 : in  unsigned(35 downto 0);
i2 : in  unsigned(35 downto 0);
i3 : in  unsigned(6 downto 0);
i4 : in  unsigned(0 downto 0);
i5 : in  unsigned(0 downto 0);
o1 : out unsigned(35 downto 0);
o2 : out unsigned(35 downto 0));
end component cf_fft_4096_18_18;
component cf_fft_4096_18_37 is
port (
clock_c : in std_logic;
i1 : in  unsigned(1 downto 0);
i2 : in  unsigned(0 downto 0);
i3 : in  unsigned(0 downto 0);
o1 : out unsigned(0 downto 0));
end component cf_fft_4096_18_37;
component cf_fft_4096_18_28 is
port (
clock_c : in std_logic;
i1 : in  unsigned(0 downto 0);
i2 : in  unsigned(0 downto 0);
i3 : in  unsigned(0 downto 0);
o1 : out unsigned(10 downto 0);
o2 : out unsigned(0 downto 0));
end component cf_fft_4096_18_28;
component cf_fft_4096_18_33 is
port (
clock_c : in std_logic;
i1 : in  unsigned(71 downto 0);
i2 : in  unsigned(0 downto 0);
i3 : in  unsigned(9 downto 0);
i4 : in  unsigned(0 downto 0);
i5 : in  unsigned(0 downto 0);
i6 : in  unsigned(0 downto 0);
o1 : out unsigned(71 downto 0));
end component cf_fft_4096_18_33;
component cf_fft_4096_18_32 is
port (
clock_c : in std_logic;
i1 : in  unsigned(71 downto 0);
i2 : in  unsigned(0 downto 0);
i3 : in  unsigned(9 downto 0);
i4 : in  unsigned(0 downto 0);
i5 : in  unsigned(0 downto 0);
i6 : in  unsigned(0 downto 0);
o1 : out unsigned(0 downto 0);
o2 : out unsigned(0 downto 0);
o3 : out unsigned(71 downto 0));
end component cf_fft_4096_18_32;
begin
n1 <= s27_1(10 downto 10) &
  s27_1(9 downto 9) &
  s27_1(8 downto 8) &
  s27_1(7 downto 7) &
  s27_1(6 downto 6) &
  s27_1(5 downto 5) &
  s27_1(4 downto 4);
n2 <= s25_1 & s25_2;
process (clock_c) begin
  if rising_edge(clock_c) then
    if i5 = "1" then
      n3 <= "0";
    elsif i4 = "1" then
      n3 <= s27_2;
    end if;
  end if;
end process;
process (clock_c) begin
  if rising_edge(clock_c) then
    if i5 = "1" then
      n4 <= "0";
    elsif i4 = "1" then
      n4 <= n3;
    end if;
  end if;
end process;
process (clock_c) begin
  if rising_edge(clock_c) then
    if i5 = "1" then
      n5 <= "0";
    elsif i4 = "1" then
      n5 <= n4;
    end if;
  end if;
end process;
process (clock_c) begin
  if rising_edge(clock_c) then
    if i5 = "1" then
      n6 <= "0";
    elsif i4 = "1" then
      n6 <= n5;
    end if;
  end if;
end process;
n7 <= s27_1(10 downto 10) &
  s27_1(9 downto 9) &
  s27_1(8 downto 8) &
  s27_1(7 downto 7) &
  s27_1(6 downto 6) &
  s27_1(5 downto 5) &
  s27_1(4 downto 4) &
  s27_1(3 downto 3) &
  s27_1(2 downto 2) &
  s27_1(1 downto 1);
process (clock_c) begin
  if rising_edge(clock_c) then
    if i5 = "1" then
      n8 <= "0000000000";
    elsif i4 = "1" then
      n8 <= n7;
    end if;
  end if;
end process;
process (clock_c) begin
  if rising_edge(clock_c) then
    if i5 = "1" then
      n9 <= "0000000000";
    elsif i4 = "1" then
      n9 <= n8;
    end if;
  end if;
end process;
process (clock_c) begin
  if rising_edge(clock_c) then
    if i5 = "1" then
      n10 <= "0000000000";
    elsif i4 = "1" then
      n10 <= n9;
    end if;
  end if;
end process;
process (clock_c) begin
  if rising_edge(clock_c) then
    if i5 = "1" then
      n11 <= "0000000000";
    elsif i4 = "1" then
      n11 <= n10;
    end if;
  end if;
end process;
n12 <= s27_1(0 downto 0);
process (clock_c) begin
  if rising_edge(clock_c) then
    if i5 = "1" then
      n13 <= "0";
    elsif i4 = "1" then
      n13 <= n12;
    end if;
  end if;
end process;
process (clock_c) begin
  if rising_edge(clock_c) then
    if i5 = "1" then
      n14 <= "0";
    elsif i4 = "1" then
      n14 <= n13;
    end if;
  end if;
end process;
process (clock_c) begin
  if rising_edge(clock_c) then
    if i5 = "1" then
      n15 <= "0";
    elsif i4 = "1" then
      n15 <= n14;
    end if;
  end if;
end process;
process (clock_c) begin
  if rising_edge(clock_c) then
    if i5 = "1" then
      n16 <= "0";
    elsif i4 = "1" then
      n16 <= n15;
    end if;
  end if;
end process;
n17 <= not n16;
n18 <= s29_2 & s29_1;
n19 <= s29_3(71 downto 71) &
  s29_3(70 downto 70) &
  s29_3(69 downto 69) &
  s29_3(68 downto 68) &
  s29_3(67 downto 67) &
  s29_3(66 downto 66) &
  s29_3(65 downto 65) &
  s29_3(64 downto 64) &
  s29_3(63 downto 63) &
  s29_3(62 downto 62) &
  s29_3(61 downto 61) &
  s29_3(60 downto 60) &
  s29_3(59 downto 59) &
  s29_3(58 downto 58) &
  s29_3(57 downto 57) &
  s29_3(56 downto 56) &
  s29_3(55 downto 55) &
  s29_3(54 downto 54) &
  s29_3(53 downto 53) &
  s29_3(52 downto 52) &
  s29_3(51 downto 51) &
  s29_3(50 downto 50) &
  s29_3(49 downto 49) &
  s29_3(48 downto 48) &
  s29_3(47 downto 47) &
  s29_3(46 downto 46) &
  s29_3(45 downto 45) &
  s29_3(44 downto 44) &
  s29_3(43 downto 43) &
  s29_3(42 downto 42) &
  s29_3(41 downto 41) &
  s29_3(40 downto 40) &
  s29_3(39 downto 39) &
  s29_3(38 downto 38) &
  s29_3(37 downto 37) &
  s29_3(36 downto 36);
n20 <= s29_3(35 downto 35) &
  s29_3(34 downto 34) &
  s29_3(33 downto 33) &
  s29_3(32 downto 32) &
  s29_3(31 downto 31) &
  s29_3(30 downto 30) &
  s29_3(29 downto 29) &
  s29_3(28 downto 28) &
  s29_3(27 downto 27) &
  s29_3(26 downto 26) &
  s29_3(25 downto 25) &
  s29_3(24 downto 24) &
  s29_3(23 downto 23) &
  s29_3(22 downto 22) &
  s29_3(21 downto 21) &
  s29_3(20 downto 20) &
  s29_3(19 downto 19) &
  s29_3(18 downto 18) &
  s29_3(17 downto 17) &
  s29_3(16 downto 16) &
  s29_3(15 downto 15) &
  s29_3(14 downto 14) &
  s29_3(13 downto 13) &
  s29_3(12 downto 12) &
  s29_3(11 downto 11) &
  s29_3(10 downto 10) &
  s29_3(9 downto 9) &
  s29_3(8 downto 8) &
  s29_3(7 downto 7) &
  s29_3(6 downto 6) &
  s29_3(5 downto 5) &
  s29_3(4 downto 4) &
  s29_3(3 downto 3) &
  s29_3(2 downto 2) &
  s29_3(1 downto 1) &
  s29_3(0 downto 0);
n21 <= s28_1(71 downto 71) &
  s28_1(70 downto 70) &
  s28_1(69 downto 69) &
  s28_1(68 downto 68) &
  s28_1(67 downto 67) &
  s28_1(66 downto 66) &
  s28_1(65 downto 65) &
  s28_1(64 downto 64) &
  s28_1(63 downto 63) &
  s28_1(62 downto 62) &
  s28_1(61 downto 61) &
  s28_1(60 downto 60) &
  s28_1(59 downto 59) &
  s28_1(58 downto 58) &
  s28_1(57 downto 57) &
  s28_1(56 downto 56) &
  s28_1(55 downto 55) &
  s28_1(54 downto 54) &
  s28_1(53 downto 53) &
  s28_1(52 downto 52) &
  s28_1(51 downto 51) &
  s28_1(50 downto 50) &
  s28_1(49 downto 49) &
  s28_1(48 downto 48) &
  s28_1(47 downto 47) &
  s28_1(46 downto 46) &
  s28_1(45 downto 45) &
  s28_1(44 downto 44) &
  s28_1(43 downto 43) &
  s28_1(42 downto 42) &
  s28_1(41 downto 41) &
  s28_1(40 downto 40) &
  s28_1(39 downto 39) &
  s28_1(38 downto 38) &
  s28_1(37 downto 37) &
  s28_1(36 downto 36);
n22 <= s28_1(35 downto 35) &
  s28_1(34 downto 34) &
  s28_1(33 downto 33) &
  s28_1(32 downto 32) &
  s28_1(31 downto 31) &
  s28_1(30 downto 30) &
  s28_1(29 downto 29) &
  s28_1(28 downto 28) &
  s28_1(27 downto 27) &
  s28_1(26 downto 26) &
  s28_1(25 downto 25) &
  s28_1(24 downto 24) &
  s28_1(23 downto 23) &
  s28_1(22 downto 22) &
  s28_1(21 downto 21) &
  s28_1(20 downto 20) &
  s28_1(19 downto 19) &
  s28_1(18 downto 18) &
  s28_1(17 downto 17) &
  s28_1(16 downto 16) &
  s28_1(15 downto 15) &
  s28_1(14 downto 14) &
  s28_1(13 downto 13) &
  s28_1(12 downto 12) &
  s28_1(11 downto 11) &
  s28_1(10 downto 10) &
  s28_1(9 downto 9) &
  s28_1(8 downto 8) &
  s28_1(7 downto 7) &
  s28_1(6 downto 6) &
  s28_1(5 downto 5) &
  s28_1(4 downto 4) &
  s28_1(3 downto 3) &
  s28_1(2 downto 2) &
  s28_1(1 downto 1) &
  s28_1(0 downto 0);
n23 <= n20 when s26_1 = "1" else n19;
n24 <= n22 when s26_1 = "1" else n21;
s25 : cf_fft_4096_18_18 port map (clock_c, i2, i3, n1, i4, i5, s25_1, s25_2);
s26 : cf_fft_4096_18_37 port map (clock_c, n18, i4, i5, s26_1);
s27 : cf_fft_4096_18_28 port map (clock_c, i1, i4, i5, s27_1, s27_2);
s28 : cf_fft_4096_18_33 port map (clock_c, n2, n6, n11, n16, i4, i5, s28_1);
s29 : cf_fft_4096_18_32 port map (clock_c, n2, n6, n11, n17, i4, i5, s29_1, s29_2, s29_3);
o3 <= n24;
o2 <= n23;
o1 <= s29_1;
end architecture rtl;

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
entity cf_fft_4096_18_16 is
port (
clock_c : in std_logic;
i1 : in  unsigned(35 downto 0);
i2 : in  unsigned(35 downto 0);
i3 : in  unsigned(5 downto 0);
i4 : in  unsigned(0 downto 0);
i5 : in  unsigned(0 downto 0);
o1 : out unsigned(35 downto 0);
o2 : out unsigned(35 downto 0));
end entity cf_fft_4096_18_16;
architecture rtl of cf_fft_4096_18_16 is
signal n1 : unsigned(35 downto 0) := "000000000000000000000000000000000000";
signal n2 : unsigned(17 downto 0);
signal n3 : unsigned(17 downto 0);
signal n4 : unsigned(35 downto 0) := "000000000000000000000000000000000000";
signal n5 : unsigned(17 downto 0);
signal n6 : unsigned(17 downto 0);
signal n7 : unsigned(17 downto 0) := "000000000000000000";
signal n8 : unsigned(17 downto 0) := "000000000000000000";
signal n9 : unsigned(17 downto 0) := "000000000000000000";
signal n10 : unsigned(17 downto 0) := "000000000000000000";
signal n11 : unsigned(35 downto 0) := "000000000000000000000000000000000000";
signal n12 : unsigned(17 downto 0);
signal n13 : unsigned(17 downto 0);
signal n14 : unsigned(35 downto 0);
signal n15 : unsigned(17 downto 0);
signal n16 : unsigned(17 downto 0) := "000000000000000000";
signal n17 : unsigned(35 downto 0);
signal n18 : unsigned(17 downto 0);
signal n19 : unsigned(17 downto 0) := "000000000000000000";
signal n20 : unsigned(17 downto 0);
signal n21 : unsigned(17 downto 0) := "000000000000000000";
signal n22 : unsigned(35 downto 0);
signal n23 : unsigned(17 downto 0);
signal n24 : unsigned(17 downto 0) := "000000000000000000";
signal n25 : unsigned(35 downto 0);
signal n26 : unsigned(17 downto 0);
signal n27 : unsigned(17 downto 0) := "000000000000000000";
signal n28 : unsigned(17 downto 0);
signal n29 : unsigned(17 downto 0) := "000000000000000000";
signal n30 : unsigned(17 downto 0);
signal n31 : unsigned(17 downto 0);
signal n32 : unsigned(35 downto 0);
signal n33 : unsigned(35 downto 0) := "000000000000000000000000000000000000";
signal n34 : unsigned(17 downto 0);
signal n35 : unsigned(17 downto 0);
signal n36 : unsigned(35 downto 0);
signal n37 : unsigned(35 downto 0) := "000000000000000000000000000000000000";
begin
process (clock_c) begin
  if rising_edge(clock_c) then
    if i5 = "1" then
      n1 <= "000000000000000000000000000000000000";
    elsif i4 = "1" then
      n1 <= i1;
    end if;
  end if;
end process;
n2 <= n1(35 downto 35) &
  n1(34 downto 34) &
  n1(33 downto 33) &
  n1(32 downto 32) &
  n1(31 downto 31) &
  n1(30 downto 30) &
  n1(29 downto 29) &
  n1(28 downto 28) &
  n1(27 downto 27) &
  n1(26 downto 26) &
  n1(25 downto 25) &
  n1(24 downto 24) &
  n1(23 downto 23) &
  n1(22 downto 22) &
  n1(21 downto 21) &
  n1(20 downto 20) &
  n1(19 downto 19) &
  n1(18 downto 18);
n3 <= n1(17 downto 17) &
  n1(16 downto 16) &
  n1(15 downto 15) &
  n1(14 downto 14) &
  n1(13 downto 13) &
  n1(12 downto 12) &
  n1(11 downto 11) &
  n1(10 downto 10) &
  n1(9 downto 9) &
  n1(8 downto 8) &
  n1(7 downto 7) &
  n1(6 downto 6) &
  n1(5 downto 5) &
  n1(4 downto 4) &
  n1(3 downto 3) &
  n1(2 downto 2) &
  n1(1 downto 1) &
  n1(0 downto 0);
process (clock_c) begin
  if rising_edge(clock_c) then
    if i5 = "1" then
      n4 <= "000000000000000000000000000000000000";
    elsif i4 = "1" then
      n4 <= i2;
    end if;
  end if;
end process;
n5 <= n4(35 downto 35) &
  n4(34 downto 34) &
  n4(33 downto 33) &
  n4(32 downto 32) &
  n4(31 downto 31) &
  n4(30 downto 30) &
  n4(29 downto 29) &
  n4(28 downto 28) &
  n4(27 downto 27) &
  n4(26 downto 26) &
  n4(25 downto 25) &
  n4(24 downto 24) &
  n4(23 downto 23) &
  n4(22 downto 22) &
  n4(21 downto 21) &
  n4(20 downto 20) &
  n4(19 downto 19) &
  n4(18 downto 18);
n6 <= n4(17 downto 17) &
  n4(16 downto 16) &
  n4(15 downto 15) &
  n4(14 downto 14) &
  n4(13 downto 13) &
  n4(12 downto 12) &
  n4(11 downto 11) &
  n4(10 downto 10) &
  n4(9 downto 9) &
  n4(8 downto 8) &
  n4(7 downto 7) &
  n4(6 downto 6) &
  n4(5 downto 5) &
  n4(4 downto 4) &
  n4(3 downto 3) &
  n4(2 downto 2) &
  n4(1 downto 1) &
  n4(0 downto 0);
process (clock_c) begin
  if rising_edge(clock_c) then
    if i5 = "1" then
      n7 <= "000000000000000000";
    elsif i4 = "1" then
      n7 <= n2;
    end if;
  end if;
end process;
process (clock_c) begin
  if rising_edge(clock_c) then
    if i5 = "1" then
      n8 <= "000000000000000000";
    elsif i4 = "1" then
      n8 <= n7;
    end if;
  end if;
end process;
process (clock_c) begin
  if rising_edge(clock_c) then
    if i5 = "1" then
      n9 <= "000000000000000000";
    elsif i4 = "1" then
      n9 <= n3;
    end if;
  end if;
end process;
process (clock_c) begin
  if rising_edge(clock_c) then
    if i5 = "1" then
      n10 <= "000000000000000000";
    elsif i4 = "1" then
      n10 <= n9;
    end if;
  end if;
end process;
process (clock_c) begin
  if rising_edge(clock_c) then 
    if i4 = "1" then
      case i3 is
        when "000000" => n11 <= "011111111111111111000000000000000000";
        when "000001" => n11 <= "011111111101100010111110011011100000";
        when "000010" => n11 <= "011111110110001000111100110111010000";
        when "000011" => n11 <= "011111101001110101111011010011011111";
        when "000100" => n11 <= "011111011000101001111001110000011101";
        when "000101" => n11 <= "011111000010100111111000001110011000";
        when "000110" => n11 <= "011110100111110100110110101101011111";
        when "000111" => n11 <= "011110001000010010110101001110000011";
        when "001000" => n11 <= "011101100100000110110011110000010000";
        when "001001" => n11 <= "011100111011010111110010010100010111";
        when "001010" => n11 <= "011100001110001011110000111010100101";
        when "001011" => n11 <= "011011011100101000101111100011000111";
        when "001100" => n11 <= "011010100110110110101110001110001100";
        when "001101" => n11 <= "011001101100111110101100111100000000";
        when "001110" => n11 <= "011000101111001000101011101100110000";
        when "001111" => n11 <= "010111101101011101101010100000101001";
        when "010000" => n11 <= "010110101000001001101001010111110110";
        when "010001" => n11 <= "010101011111010110101000010010100010";
        when "010010" => n11 <= "010100010011001111100111010000110111";
        when "010011" => n11 <= "010011000011111111100110010011000001";
        when "010100" => n11 <= "010001110001110011100101011001001001";
        when "010101" => n11 <= "010000011100111000100100100011010111";
        when "010110" => n11 <= "001111000101011010100011110001110100";
        when "010111" => n11 <= "001101101011101000100011000100101000";
        when "011000" => n11 <= "001100001111101111100010011011111001";
        when "011001" => n11 <= "001010110001111100100001110111101101";
        when "011010" => n11 <= "001001010010100000100001011000001011";
        when "011011" => n11 <= "000111110001100111100000111101011000";
        when "011100" => n11 <= "000110001111100010100000100111010110";
        when "011101" => n11 <= "000100101100100000100000010110001010";
        when "011110" => n11 <= "000011001000101111100000001001110111";
        when "011111" => n11 <= "000001100100011111100000000010011101";
        when "100000" => n11 <= "000000000000000000100000000000000000";
        when "100001" => n11 <= "111110011011100000100000000010011101";
        when "100010" => n11 <= "111100110111010000100000001001110111";
        when "100011" => n11 <= "111011010011011111100000010110001010";
        when "100100" => n11 <= "111001110000011101100000100111010110";
        when "100101" => n11 <= "111000001110011000100000111101011000";
        when "100110" => n11 <= "110110101101011111100001011000001011";
        when "100111" => n11 <= "110101001110000011100001110111101101";
        when "101000" => n11 <= "110011110000010000100010011011111001";
        when "101001" => n11 <= "110010010100010111100011000100101000";
        when "101010" => n11 <= "110000111010100101100011110001110100";
        when "101011" => n11 <= "101111100011000111100100100011010111";
        when "101100" => n11 <= "101110001110001100100101011001001001";
        when "101101" => n11 <= "101100111100000000100110010011000001";
        when "101110" => n11 <= "101011101100110000100111010000110111";
        when "101111" => n11 <= "101010100000101001101000010010100010";
        when "110000" => n11 <= "101001010111110110101001010111110110";
        when "110001" => n11 <= "101000010010100010101010100000101001";
        when "110010" => n11 <= "100111010000110111101011101100110000";
        when "110011" => n11 <= "100110010011000001101100111100000000";
        when "110100" => n11 <= "100101011001001001101110001110001100";
        when "110101" => n11 <= "100100100011010111101111100011000111";
        when "110110" => n11 <= "100011110001110100110000111010100101";
        when "110111" => n11 <= "100011000100101000110010010100010111";
        when "111000" => n11 <= "100010011011111001110011110000010000";
        when "111001" => n11 <= "100001110111101101110101001110000011";
        when "111010" => n11 <= "100001011000001011110110101101011111";
        when "111011" => n11 <= "100000111101011000111000001110011000";
        when "111100" => n11 <= "100000100111010110111001110000011101";
        when "111101" => n11 <= "100000010110001010111011010011011111";
        when "111110" => n11 <= "100000001001110111111100110111010000";
        when "111111" => n11 <= "100000000010011101111110011011100000";
        when others => n11 <= "XXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX";
      end case;
    end if;
  end if;
end process;
n12 <= n11(35 downto 35) &
  n11(34 downto 34) &
  n11(33 downto 33) &
  n11(32 downto 32) &
  n11(31 downto 31) &
  n11(30 downto 30) &
  n11(29 downto 29) &
  n11(28 downto 28) &
  n11(27 downto 27) &
  n11(26 downto 26) &
  n11(25 downto 25) &
  n11(24 downto 24) &
  n11(23 downto 23) &
  n11(22 downto 22) &
  n11(21 downto 21) &
  n11(20 downto 20) &
  n11(19 downto 19) &
  n11(18 downto 18);
n13 <= n11(17 downto 17) &
  n11(16 downto 16) &
  n11(15 downto 15) &
  n11(14 downto 14) &
  n11(13 downto 13) &
  n11(12 downto 12) &
  n11(11 downto 11) &
  n11(10 downto 10) &
  n11(9 downto 9) &
  n11(8 downto 8) &
  n11(7 downto 7) &
  n11(6 downto 6) &
  n11(5 downto 5) &
  n11(4 downto 4) &
  n11(3 downto 3) &
  n11(2 downto 2) &
  n11(1 downto 1) &
  n11(0 downto 0);
n14 <= unsigned(signed(n5) * signed(n12));
n15 <= n14(34 downto 34) &
  n14(33 downto 33) &
  n14(32 downto 32) &
  n14(31 downto 31) &
  n14(30 downto 30) &
  n14(29 downto 29) &
  n14(28 downto 28) &
  n14(27 downto 27) &
  n14(26 downto 26) &
  n14(25 downto 25) &
  n14(24 downto 24) &
  n14(23 downto 23) &
  n14(22 downto 22) &
  n14(21 downto 21) &
  n14(20 downto 20) &
  n14(19 downto 19) &
  n14(18 downto 18) &
  n14(17 downto 17);
process (clock_c) begin
  if rising_edge(clock_c) then
    if i5 = "1" then
      n16 <= "000000000000000000";
    elsif i4 = "1" then
      n16 <= n15;
    end if;
  end if;
end process;
n17 <= unsigned(signed(n6) * signed(n13));
n18 <= n17(34 downto 34) &
  n17(33 downto 33) &
  n17(32 downto 32) &
  n17(31 downto 31) &
  n17(30 downto 30) &
  n17(29 downto 29) &
  n17(28 downto 28) &
  n17(27 downto 27) &
  n17(26 downto 26) &
  n17(25 downto 25) &
  n17(24 downto 24) &
  n17(23 downto 23) &
  n17(22 downto 22) &
  n17(21 downto 21) &
  n17(20 downto 20) &
  n17(19 downto 19) &
  n17(18 downto 18) &
  n17(17 downto 17);
process (clock_c) begin
  if rising_edge(clock_c) then
    if i5 = "1" then
      n19 <= "000000000000000000";
    elsif i4 = "1" then
      n19 <= n18;
    end if;
  end if;
end process;
n20 <= n16 - n19;
process (clock_c) begin
  if rising_edge(clock_c) then
    if i5 = "1" then
      n21 <= "000000000000000000";
    elsif i4 = "1" then
      n21 <= n20;
    end if;
  end if;
end process;
n22 <= unsigned(signed(n5) * signed(n13));
n23 <= n22(34 downto 34) &
  n22(33 downto 33) &
  n22(32 downto 32) &
  n22(31 downto 31) &
  n22(30 downto 30) &
  n22(29 downto 29) &
  n22(28 downto 28) &
  n22(27 downto 27) &
  n22(26 downto 26) &
  n22(25 downto 25) &
  n22(24 downto 24) &
  n22(23 downto 23) &
  n22(22 downto 22) &
  n22(21 downto 21) &
  n22(20 downto 20) &
  n22(19 downto 19) &
  n22(18 downto 18) &
  n22(17 downto 17);
process (clock_c) begin
  if rising_edge(clock_c) then
    if i5 = "1" then
      n24 <= "000000000000000000";
    elsif i4 = "1" then
      n24 <= n23;
    end if;
  end if;
end process;
n25 <= unsigned(signed(n6) * signed(n12));
n26 <= n25(34 downto 34) &
  n25(33 downto 33) &
  n25(32 downto 32) &
  n25(31 downto 31) &
  n25(30 downto 30) &
  n25(29 downto 29) &
  n25(28 downto 28) &
  n25(27 downto 27) &
  n25(26 downto 26) &
  n25(25 downto 25) &
  n25(24 downto 24) &
  n25(23 downto 23) &
  n25(22 downto 22) &
  n25(21 downto 21) &
  n25(20 downto 20) &
  n25(19 downto 19) &
  n25(18 downto 18) &
  n25(17 downto 17);
process (clock_c) begin
  if rising_edge(clock_c) then
    if i5 = "1" then
      n27 <= "000000000000000000";
    elsif i4 = "1" then
      n27 <= n26;
    end if;
  end if;
end process;
n28 <= n24 + n27;
process (clock_c) begin
  if rising_edge(clock_c) then
    if i5 = "1" then
      n29 <= "000000000000000000";
    elsif i4 = "1" then
      n29 <= n28;
    end if;
  end if;
end process;
n30 <= n8 + n21;
n31 <= n10 + n29;
n32 <= n30 & n31;
process (clock_c) begin
  if rising_edge(clock_c) then
    if i5 = "1" then
      n33 <= "000000000000000000000000000000000000";
    elsif i4 = "1" then
      n33 <= n32;
    end if;
  end if;
end process;
n34 <= n8 - n21;
n35 <= n10 - n29;
n36 <= n34 & n35;
process (clock_c) begin
  if rising_edge(clock_c) then
    if i5 = "1" then
      n37 <= "000000000000000000000000000000000000";
    elsif i4 = "1" then
      n37 <= n36;
    end if;
  end if;
end process;
o2 <= n37;
o1 <= n33;
end architecture rtl;

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
entity cf_fft_4096_18_15 is
port (
clock_c : in std_logic;
i1 : in  unsigned(0 downto 0);
i2 : in  unsigned(35 downto 0);
i3 : in  unsigned(35 downto 0);
i4 : in  unsigned(0 downto 0);
i5 : in  unsigned(0 downto 0);
o1 : out unsigned(0 downto 0);
o2 : out unsigned(35 downto 0);
o3 : out unsigned(35 downto 0));
end entity cf_fft_4096_18_15;
architecture rtl of cf_fft_4096_18_15 is
signal n1 : unsigned(5 downto 0);
signal n2 : unsigned(71 downto 0);
signal n3 : unsigned(0 downto 0) := "0";
signal n4 : unsigned(0 downto 0) := "0";
signal n5 : unsigned(0 downto 0) := "0";
signal n6 : unsigned(0 downto 0) := "0";
signal n7 : unsigned(9 downto 0);
signal n8 : unsigned(9 downto 0) := "0000000000";
signal n9 : unsigned(9 downto 0) := "0000000000";
signal n10 : unsigned(9 downto 0) := "0000000000";
signal n11 : unsigned(9 downto 0) := "0000000000";
signal n12 : unsigned(0 downto 0);
signal n13 : unsigned(0 downto 0) := "0";
signal n14 : unsigned(0 downto 0) := "0";
signal n15 : unsigned(0 downto 0) := "0";
signal n16 : unsigned(0 downto 0) := "0";
signal n17 : unsigned(0 downto 0);
signal n18 : unsigned(1 downto 0);
signal n19 : unsigned(35 downto 0);
signal n20 : unsigned(35 downto 0);
signal n21 : unsigned(35 downto 0);
signal n22 : unsigned(35 downto 0);
signal n23 : unsigned(35 downto 0);
signal n24 : unsigned(35 downto 0);
signal s25_1 : unsigned(0 downto 0);
signal s26_1 : unsigned(35 downto 0);
signal s26_2 : unsigned(35 downto 0);
signal s27_1 : unsigned(10 downto 0);
signal s27_2 : unsigned(0 downto 0);
signal s28_1 : unsigned(0 downto 0);
signal s28_2 : unsigned(0 downto 0);
signal s28_3 : unsigned(71 downto 0);
signal s29_1 : unsigned(71 downto 0);
component cf_fft_4096_18_37 is
port (
clock_c : in std_logic;
i1 : in  unsigned(1 downto 0);
i2 : in  unsigned(0 downto 0);
i3 : in  unsigned(0 downto 0);
o1 : out unsigned(0 downto 0));
end component cf_fft_4096_18_37;
component cf_fft_4096_18_16 is
port (
clock_c : in std_logic;
i1 : in  unsigned(35 downto 0);
i2 : in  unsigned(35 downto 0);
i3 : in  unsigned(5 downto 0);
i4 : in  unsigned(0 downto 0);
i5 : in  unsigned(0 downto 0);
o1 : out unsigned(35 downto 0);
o2 : out unsigned(35 downto 0));
end component cf_fft_4096_18_16;
component cf_fft_4096_18_28 is
port (
clock_c : in std_logic;
i1 : in  unsigned(0 downto 0);
i2 : in  unsigned(0 downto 0);
i3 : in  unsigned(0 downto 0);
o1 : out unsigned(10 downto 0);
o2 : out unsigned(0 downto 0));
end component cf_fft_4096_18_28;
component cf_fft_4096_18_32 is
port (
clock_c : in std_logic;
i1 : in  unsigned(71 downto 0);
i2 : in  unsigned(0 downto 0);
i3 : in  unsigned(9 downto 0);
i4 : in  unsigned(0 downto 0);
i5 : in  unsigned(0 downto 0);
i6 : in  unsigned(0 downto 0);
o1 : out unsigned(0 downto 0);
o2 : out unsigned(0 downto 0);
o3 : out unsigned(71 downto 0));
end component cf_fft_4096_18_32;
component cf_fft_4096_18_33 is
port (
clock_c : in std_logic;
i1 : in  unsigned(71 downto 0);
i2 : in  unsigned(0 downto 0);
i3 : in  unsigned(9 downto 0);
i4 : in  unsigned(0 downto 0);
i5 : in  unsigned(0 downto 0);
i6 : in  unsigned(0 downto 0);
o1 : out unsigned(71 downto 0));
end component cf_fft_4096_18_33;
begin
n1 <= s27_1(10 downto 10) &
  s27_1(9 downto 9) &
  s27_1(8 downto 8) &
  s27_1(7 downto 7) &
  s27_1(6 downto 6) &
  s27_1(5 downto 5);
n2 <= s26_1 & s26_2;
process (clock_c) begin
  if rising_edge(clock_c) then
    if i5 = "1" then
      n3 <= "0";
    elsif i4 = "1" then
      n3 <= s27_2;
    end if;
  end if;
end process;
process (clock_c) begin
  if rising_edge(clock_c) then
    if i5 = "1" then
      n4 <= "0";
    elsif i4 = "1" then
      n4 <= n3;
    end if;
  end if;
end process;
process (clock_c) begin
  if rising_edge(clock_c) then
    if i5 = "1" then
      n5 <= "0";
    elsif i4 = "1" then
      n5 <= n4;
    end if;
  end if;
end process;
process (clock_c) begin
  if rising_edge(clock_c) then
    if i5 = "1" then
      n6 <= "0";
    elsif i4 = "1" then
      n6 <= n5;
    end if;
  end if;
end process;
n7 <= s27_1(10 downto 10) &
  s27_1(9 downto 9) &
  s27_1(8 downto 8) &
  s27_1(7 downto 7) &
  s27_1(6 downto 6) &
  s27_1(5 downto 5) &
  s27_1(4 downto 4) &
  s27_1(3 downto 3) &
  s27_1(2 downto 2) &
  s27_1(1 downto 1);
process (clock_c) begin
  if rising_edge(clock_c) then
    if i5 = "1" then
      n8 <= "0000000000";
    elsif i4 = "1" then
      n8 <= n7;
    end if;
  end if;
end process;
process (clock_c) begin
  if rising_edge(clock_c) then
    if i5 = "1" then
      n9 <= "0000000000";
    elsif i4 = "1" then
      n9 <= n8;
    end if;
  end if;
end process;
process (clock_c) begin
  if rising_edge(clock_c) then
    if i5 = "1" then
      n10 <= "0000000000";
    elsif i4 = "1" then
      n10 <= n9;
    end if;
  end if;
end process;
process (clock_c) begin
  if rising_edge(clock_c) then
    if i5 = "1" then
      n11 <= "0000000000";
    elsif i4 = "1" then
      n11 <= n10;
    end if;
  end if;
end process;
n12 <= s27_1(0 downto 0);
process (clock_c) begin
  if rising_edge(clock_c) then
    if i5 = "1" then
      n13 <= "0";
    elsif i4 = "1" then
      n13 <= n12;
    end if;
  end if;
end process;
process (clock_c) begin
  if rising_edge(clock_c) then
    if i5 = "1" then
      n14 <= "0";
    elsif i4 = "1" then
      n14 <= n13;
    end if;
  end if;
end process;
process (clock_c) begin
  if rising_edge(clock_c) then
    if i5 = "1" then
      n15 <= "0";
    elsif i4 = "1" then
      n15 <= n14;
    end if;
  end if;
end process;
process (clock_c) begin
  if rising_edge(clock_c) then
    if i5 = "1" then
      n16 <= "0";
    elsif i4 = "1" then
      n16 <= n15;
    end if;
  end if;
end process;
n17 <= not n16;
n18 <= s28_2 & s28_1;
n19 <= s28_3(71 downto 71) &
  s28_3(70 downto 70) &
  s28_3(69 downto 69) &
  s28_3(68 downto 68) &
  s28_3(67 downto 67) &
  s28_3(66 downto 66) &
  s28_3(65 downto 65) &
  s28_3(64 downto 64) &
  s28_3(63 downto 63) &
  s28_3(62 downto 62) &
  s28_3(61 downto 61) &
  s28_3(60 downto 60) &
  s28_3(59 downto 59) &
  s28_3(58 downto 58) &
  s28_3(57 downto 57) &
  s28_3(56 downto 56) &
  s28_3(55 downto 55) &
  s28_3(54 downto 54) &
  s28_3(53 downto 53) &
  s28_3(52 downto 52) &
  s28_3(51 downto 51) &
  s28_3(50 downto 50) &
  s28_3(49 downto 49) &
  s28_3(48 downto 48) &
  s28_3(47 downto 47) &
  s28_3(46 downto 46) &
  s28_3(45 downto 45) &
  s28_3(44 downto 44) &
  s28_3(43 downto 43) &
  s28_3(42 downto 42) &
  s28_3(41 downto 41) &
  s28_3(40 downto 40) &
  s28_3(39 downto 39) &
  s28_3(38 downto 38) &
  s28_3(37 downto 37) &
  s28_3(36 downto 36);
n20 <= s28_3(35 downto 35) &
  s28_3(34 downto 34) &
  s28_3(33 downto 33) &
  s28_3(32 downto 32) &
  s28_3(31 downto 31) &
  s28_3(30 downto 30) &
  s28_3(29 downto 29) &
  s28_3(28 downto 28) &
  s28_3(27 downto 27) &
  s28_3(26 downto 26) &
  s28_3(25 downto 25) &
  s28_3(24 downto 24) &
  s28_3(23 downto 23) &
  s28_3(22 downto 22) &
  s28_3(21 downto 21) &
  s28_3(20 downto 20) &
  s28_3(19 downto 19) &
  s28_3(18 downto 18) &
  s28_3(17 downto 17) &
  s28_3(16 downto 16) &
  s28_3(15 downto 15) &
  s28_3(14 downto 14) &
  s28_3(13 downto 13) &
  s28_3(12 downto 12) &
  s28_3(11 downto 11) &
  s28_3(10 downto 10) &
  s28_3(9 downto 9) &
  s28_3(8 downto 8) &
  s28_3(7 downto 7) &
  s28_3(6 downto 6) &
  s28_3(5 downto 5) &
  s28_3(4 downto 4) &
  s28_3(3 downto 3) &
  s28_3(2 downto 2) &
  s28_3(1 downto 1) &
  s28_3(0 downto 0);
n21 <= s29_1(71 downto 71) &
  s29_1(70 downto 70) &
  s29_1(69 downto 69) &
  s29_1(68 downto 68) &
  s29_1(67 downto 67) &
  s29_1(66 downto 66) &
  s29_1(65 downto 65) &
  s29_1(64 downto 64) &
  s29_1(63 downto 63) &
  s29_1(62 downto 62) &
  s29_1(61 downto 61) &
  s29_1(60 downto 60) &
  s29_1(59 downto 59) &
  s29_1(58 downto 58) &
  s29_1(57 downto 57) &
  s29_1(56 downto 56) &
  s29_1(55 downto 55) &
  s29_1(54 downto 54) &
  s29_1(53 downto 53) &
  s29_1(52 downto 52) &
  s29_1(51 downto 51) &
  s29_1(50 downto 50) &
  s29_1(49 downto 49) &
  s29_1(48 downto 48) &
  s29_1(47 downto 47) &
  s29_1(46 downto 46) &
  s29_1(45 downto 45) &
  s29_1(44 downto 44) &
  s29_1(43 downto 43) &
  s29_1(42 downto 42) &
  s29_1(41 downto 41) &
  s29_1(40 downto 40) &
  s29_1(39 downto 39) &
  s29_1(38 downto 38) &
  s29_1(37 downto 37) &
  s29_1(36 downto 36);
n22 <= s29_1(35 downto 35) &
  s29_1(34 downto 34) &
  s29_1(33 downto 33) &
  s29_1(32 downto 32) &
  s29_1(31 downto 31) &
  s29_1(30 downto 30) &
  s29_1(29 downto 29) &
  s29_1(28 downto 28) &
  s29_1(27 downto 27) &
  s29_1(26 downto 26) &
  s29_1(25 downto 25) &
  s29_1(24 downto 24) &
  s29_1(23 downto 23) &
  s29_1(22 downto 22) &
  s29_1(21 downto 21) &
  s29_1(20 downto 20) &
  s29_1(19 downto 19) &
  s29_1(18 downto 18) &
  s29_1(17 downto 17) &
  s29_1(16 downto 16) &
  s29_1(15 downto 15) &
  s29_1(14 downto 14) &
  s29_1(13 downto 13) &
  s29_1(12 downto 12) &
  s29_1(11 downto 11) &
  s29_1(10 downto 10) &
  s29_1(9 downto 9) &
  s29_1(8 downto 8) &
  s29_1(7 downto 7) &
  s29_1(6 downto 6) &
  s29_1(5 downto 5) &
  s29_1(4 downto 4) &
  s29_1(3 downto 3) &
  s29_1(2 downto 2) &
  s29_1(1 downto 1) &
  s29_1(0 downto 0);
n23 <= n20 when s25_1 = "1" else n19;
n24 <= n22 when s25_1 = "1" else n21;
s25 : cf_fft_4096_18_37 port map (clock_c, n18, i4, i5, s25_1);
s26 : cf_fft_4096_18_16 port map (clock_c, i2, i3, n1, i4, i5, s26_1, s26_2);
s27 : cf_fft_4096_18_28 port map (clock_c, i1, i4, i5, s27_1, s27_2);
s28 : cf_fft_4096_18_32 port map (clock_c, n2, n6, n11, n17, i4, i5, s28_1, s28_2, s28_3);
s29 : cf_fft_4096_18_33 port map (clock_c, n2, n6, n11, n16, i4, i5, s29_1);
o3 <= n24;
o2 <= n23;
o1 <= s28_1;
end architecture rtl;

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
entity cf_fft_4096_18_14 is
port (
clock_c : in std_logic;
i1 : in  unsigned(35 downto 0);
i2 : in  unsigned(35 downto 0);
i3 : in  unsigned(4 downto 0);
i4 : in  unsigned(0 downto 0);
i5 : in  unsigned(0 downto 0);
o1 : out unsigned(35 downto 0);
o2 : out unsigned(35 downto 0));
end entity cf_fft_4096_18_14;
architecture rtl of cf_fft_4096_18_14 is
signal n1 : unsigned(35 downto 0) := "000000000000000000000000000000000000";
signal n2 : unsigned(17 downto 0);
signal n3 : unsigned(17 downto 0);
signal n4 : unsigned(35 downto 0) := "000000000000000000000000000000000000";
signal n5 : unsigned(17 downto 0);
signal n6 : unsigned(17 downto 0);
signal n7 : unsigned(17 downto 0) := "000000000000000000";
signal n8 : unsigned(17 downto 0) := "000000000000000000";
signal n9 : unsigned(17 downto 0) := "000000000000000000";
signal n10 : unsigned(17 downto 0) := "000000000000000000";
signal n11 : unsigned(35 downto 0) := "000000000000000000000000000000000000";
signal n12 : unsigned(17 downto 0);
signal n13 : unsigned(17 downto 0);
signal n14 : unsigned(35 downto 0);
signal n15 : unsigned(17 downto 0);
signal n16 : unsigned(17 downto 0) := "000000000000000000";
signal n17 : unsigned(35 downto 0);
signal n18 : unsigned(17 downto 0);
signal n19 : unsigned(17 downto 0) := "000000000000000000";
signal n20 : unsigned(17 downto 0);
signal n21 : unsigned(17 downto 0) := "000000000000000000";
signal n22 : unsigned(35 downto 0);
signal n23 : unsigned(17 downto 0);
signal n24 : unsigned(17 downto 0) := "000000000000000000";
signal n25 : unsigned(35 downto 0);
signal n26 : unsigned(17 downto 0);
signal n27 : unsigned(17 downto 0) := "000000000000000000";
signal n28 : unsigned(17 downto 0);
signal n29 : unsigned(17 downto 0) := "000000000000000000";
signal n30 : unsigned(17 downto 0);
signal n31 : unsigned(17 downto 0);
signal n32 : unsigned(35 downto 0);
signal n33 : unsigned(35 downto 0) := "000000000000000000000000000000000000";
signal n34 : unsigned(17 downto 0);
signal n35 : unsigned(17 downto 0);
signal n36 : unsigned(35 downto 0);
signal n37 : unsigned(35 downto 0) := "000000000000000000000000000000000000";
begin
process (clock_c) begin
  if rising_edge(clock_c) then
    if i5 = "1" then
      n1 <= "000000000000000000000000000000000000";
    elsif i4 = "1" then
      n1 <= i1;
    end if;
  end if;
end process;
n2 <= n1(35 downto 35) &
  n1(34 downto 34) &
  n1(33 downto 33) &
  n1(32 downto 32) &
  n1(31 downto 31) &
  n1(30 downto 30) &
  n1(29 downto 29) &
  n1(28 downto 28) &
  n1(27 downto 27) &
  n1(26 downto 26) &
  n1(25 downto 25) &
  n1(24 downto 24) &
  n1(23 downto 23) &
  n1(22 downto 22) &
  n1(21 downto 21) &
  n1(20 downto 20) &
  n1(19 downto 19) &
  n1(18 downto 18);
n3 <= n1(17 downto 17) &
  n1(16 downto 16) &
  n1(15 downto 15) &
  n1(14 downto 14) &
  n1(13 downto 13) &
  n1(12 downto 12) &
  n1(11 downto 11) &
  n1(10 downto 10) &
  n1(9 downto 9) &
  n1(8 downto 8) &
  n1(7 downto 7) &
  n1(6 downto 6) &
  n1(5 downto 5) &
  n1(4 downto 4) &
  n1(3 downto 3) &
  n1(2 downto 2) &
  n1(1 downto 1) &
  n1(0 downto 0);
process (clock_c) begin
  if rising_edge(clock_c) then
    if i5 = "1" then
      n4 <= "000000000000000000000000000000000000";
    elsif i4 = "1" then
      n4 <= i2;
    end if;
  end if;
end process;
n5 <= n4(35 downto 35) &
  n4(34 downto 34) &
  n4(33 downto 33) &
  n4(32 downto 32) &
  n4(31 downto 31) &
  n4(30 downto 30) &
  n4(29 downto 29) &
  n4(28 downto 28) &
  n4(27 downto 27) &
  n4(26 downto 26) &
  n4(25 downto 25) &
  n4(24 downto 24) &
  n4(23 downto 23) &
  n4(22 downto 22) &
  n4(21 downto 21) &
  n4(20 downto 20) &
  n4(19 downto 19) &
  n4(18 downto 18);
n6 <= n4(17 downto 17) &
  n4(16 downto 16) &
  n4(15 downto 15) &
  n4(14 downto 14) &
  n4(13 downto 13) &
  n4(12 downto 12) &
  n4(11 downto 11) &
  n4(10 downto 10) &
  n4(9 downto 9) &
  n4(8 downto 8) &
  n4(7 downto 7) &
  n4(6 downto 6) &
  n4(5 downto 5) &
  n4(4 downto 4) &
  n4(3 downto 3) &
  n4(2 downto 2) &
  n4(1 downto 1) &
  n4(0 downto 0);
process (clock_c) begin
  if rising_edge(clock_c) then
    if i5 = "1" then
      n7 <= "000000000000000000";
    elsif i4 = "1" then
      n7 <= n2;
    end if;
  end if;
end process;
process (clock_c) begin
  if rising_edge(clock_c) then
    if i5 = "1" then
      n8 <= "000000000000000000";
    elsif i4 = "1" then
      n8 <= n7;
    end if;
  end if;
end process;
process (clock_c) begin
  if rising_edge(clock_c) then
    if i5 = "1" then
      n9 <= "000000000000000000";
    elsif i4 = "1" then
      n9 <= n3;
    end if;
  end if;
end process;
process (clock_c) begin
  if rising_edge(clock_c) then
    if i5 = "1" then
      n10 <= "000000000000000000";
    elsif i4 = "1" then
      n10 <= n9;
    end if;
  end if;
end process;
process (clock_c) begin
  if rising_edge(clock_c) then 
    if i4 = "1" then
      case i3 is
        when "00000" => n11 <= "011111111111111111000000000000000000";
        when "00001" => n11 <= "011111110110001000111100110111010000";
        when "00010" => n11 <= "011111011000101001111001110000011101";
        when "00011" => n11 <= "011110100111110100110110101101011111";
        when "00100" => n11 <= "011101100100000110110011110000010000";
        when "00101" => n11 <= "011100001110001011110000111010100101";
        when "00110" => n11 <= "011010100110110110101110001110001100";
        when "00111" => n11 <= "011000101111001000101011101100110000";
        when "01000" => n11 <= "010110101000001001101001010111110110";
        when "01001" => n11 <= "010100010011001111100111010000110111";
        when "01010" => n11 <= "010001110001110011100101011001001001";
        when "01011" => n11 <= "001111000101011010100011110001110100";
        when "01100" => n11 <= "001100001111101111100010011011111001";
        when "01101" => n11 <= "001001010010100000100001011000001011";
        when "01110" => n11 <= "000110001111100010100000100111010110";
        when "01111" => n11 <= "000011001000101111100000001001110111";
        when "10000" => n11 <= "000000000000000000100000000000000000";
        when "10001" => n11 <= "111100110111010000100000001001110111";
        when "10010" => n11 <= "111001110000011101100000100111010110";
        when "10011" => n11 <= "110110101101011111100001011000001011";
        when "10100" => n11 <= "110011110000010000100010011011111001";
        when "10101" => n11 <= "110000111010100101100011110001110100";
        when "10110" => n11 <= "101110001110001100100101011001001001";
        when "10111" => n11 <= "101011101100110000100111010000110111";
        when "11000" => n11 <= "101001010111110110101001010111110110";
        when "11001" => n11 <= "100111010000110111101011101100110000";
        when "11010" => n11 <= "100101011001001001101110001110001100";
        when "11011" => n11 <= "100011110001110100110000111010100101";
        when "11100" => n11 <= "100010011011111001110011110000010000";
        when "11101" => n11 <= "100001011000001011110110101101011111";
        when "11110" => n11 <= "100000100111010110111001110000011101";
        when "11111" => n11 <= "100000001001110111111100110111010000";
        when others => n11 <= "XXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX";
      end case;
    end if;
  end if;
end process;
n12 <= n11(35 downto 35) &
  n11(34 downto 34) &
  n11(33 downto 33) &
  n11(32 downto 32) &
  n11(31 downto 31) &
  n11(30 downto 30) &
  n11(29 downto 29) &
  n11(28 downto 28) &
  n11(27 downto 27) &
  n11(26 downto 26) &
  n11(25 downto 25) &
  n11(24 downto 24) &
  n11(23 downto 23) &
  n11(22 downto 22) &
  n11(21 downto 21) &
  n11(20 downto 20) &
  n11(19 downto 19) &
  n11(18 downto 18);
n13 <= n11(17 downto 17) &
  n11(16 downto 16) &
  n11(15 downto 15) &
  n11(14 downto 14) &
  n11(13 downto 13) &
  n11(12 downto 12) &
  n11(11 downto 11) &
  n11(10 downto 10) &
  n11(9 downto 9) &
  n11(8 downto 8) &
  n11(7 downto 7) &
  n11(6 downto 6) &
  n11(5 downto 5) &
  n11(4 downto 4) &
  n11(3 downto 3) &
  n11(2 downto 2) &
  n11(1 downto 1) &
  n11(0 downto 0);
n14 <= unsigned(signed(n5) * signed(n12));
n15 <= n14(34 downto 34) &
  n14(33 downto 33) &
  n14(32 downto 32) &
  n14(31 downto 31) &
  n14(30 downto 30) &
  n14(29 downto 29) &
  n14(28 downto 28) &
  n14(27 downto 27) &
  n14(26 downto 26) &
  n14(25 downto 25) &
  n14(24 downto 24) &
  n14(23 downto 23) &
  n14(22 downto 22) &
  n14(21 downto 21) &
  n14(20 downto 20) &
  n14(19 downto 19) &
  n14(18 downto 18) &
  n14(17 downto 17);
process (clock_c) begin
  if rising_edge(clock_c) then
    if i5 = "1" then
      n16 <= "000000000000000000";
    elsif i4 = "1" then
      n16 <= n15;
    end if;
  end if;
end process;
n17 <= unsigned(signed(n6) * signed(n13));
n18 <= n17(34 downto 34) &
  n17(33 downto 33) &
  n17(32 downto 32) &
  n17(31 downto 31) &
  n17(30 downto 30) &
  n17(29 downto 29) &
  n17(28 downto 28) &
  n17(27 downto 27) &
  n17(26 downto 26) &
  n17(25 downto 25) &
  n17(24 downto 24) &
  n17(23 downto 23) &
  n17(22 downto 22) &
  n17(21 downto 21) &
  n17(20 downto 20) &
  n17(19 downto 19) &
  n17(18 downto 18) &
  n17(17 downto 17);
process (clock_c) begin
  if rising_edge(clock_c) then
    if i5 = "1" then
      n19 <= "000000000000000000";
    elsif i4 = "1" then
      n19 <= n18;
    end if;
  end if;
end process;
n20 <= n16 - n19;
process (clock_c) begin
  if rising_edge(clock_c) then
    if i5 = "1" then
      n21 <= "000000000000000000";
    elsif i4 = "1" then
      n21 <= n20;
    end if;
  end if;
end process;
n22 <= unsigned(signed(n5) * signed(n13));
n23 <= n22(34 downto 34) &
  n22(33 downto 33) &
  n22(32 downto 32) &
  n22(31 downto 31) &
  n22(30 downto 30) &
  n22(29 downto 29) &
  n22(28 downto 28) &
  n22(27 downto 27) &
  n22(26 downto 26) &
  n22(25 downto 25) &
  n22(24 downto 24) &
  n22(23 downto 23) &
  n22(22 downto 22) &
  n22(21 downto 21) &
  n22(20 downto 20) &
  n22(19 downto 19) &
  n22(18 downto 18) &
  n22(17 downto 17);
process (clock_c) begin
  if rising_edge(clock_c) then
    if i5 = "1" then
      n24 <= "000000000000000000";
    elsif i4 = "1" then
      n24 <= n23;
    end if;
  end if;
end process;
n25 <= unsigned(signed(n6) * signed(n12));
n26 <= n25(34 downto 34) &
  n25(33 downto 33) &
  n25(32 downto 32) &
  n25(31 downto 31) &
  n25(30 downto 30) &
  n25(29 downto 29) &
  n25(28 downto 28) &
  n25(27 downto 27) &
  n25(26 downto 26) &
  n25(25 downto 25) &
  n25(24 downto 24) &
  n25(23 downto 23) &
  n25(22 downto 22) &
  n25(21 downto 21) &
  n25(20 downto 20) &
  n25(19 downto 19) &
  n25(18 downto 18) &
  n25(17 downto 17);
process (clock_c) begin
  if rising_edge(clock_c) then
    if i5 = "1" then
      n27 <= "000000000000000000";
    elsif i4 = "1" then
      n27 <= n26;
    end if;
  end if;
end process;
n28 <= n24 + n27;
process (clock_c) begin
  if rising_edge(clock_c) then
    if i5 = "1" then
      n29 <= "000000000000000000";
    elsif i4 = "1" then
      n29 <= n28;
    end if;
  end if;
end process;
n30 <= n8 + n21;
n31 <= n10 + n29;
n32 <= n30 & n31;
process (clock_c) begin
  if rising_edge(clock_c) then
    if i5 = "1" then
      n33 <= "000000000000000000000000000000000000";
    elsif i4 = "1" then
      n33 <= n32;
    end if;
  end if;
end process;
n34 <= n8 - n21;
n35 <= n10 - n29;
n36 <= n34 & n35;
process (clock_c) begin
  if rising_edge(clock_c) then
    if i5 = "1" then
      n37 <= "000000000000000000000000000000000000";
    elsif i4 = "1" then
      n37 <= n36;
    end if;
  end if;
end process;
o2 <= n37;
o1 <= n33;
end architecture rtl;

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
entity cf_fft_4096_18_13 is
port (
clock_c : in std_logic;
i1 : in  unsigned(0 downto 0);
i2 : in  unsigned(35 downto 0);
i3 : in  unsigned(35 downto 0);
i4 : in  unsigned(0 downto 0);
i5 : in  unsigned(0 downto 0);
o1 : out unsigned(0 downto 0);
o2 : out unsigned(35 downto 0);
o3 : out unsigned(35 downto 0));
end entity cf_fft_4096_18_13;
architecture rtl of cf_fft_4096_18_13 is
signal n1 : unsigned(4 downto 0);
signal n2 : unsigned(71 downto 0);
signal n3 : unsigned(0 downto 0) := "0";
signal n4 : unsigned(0 downto 0) := "0";
signal n5 : unsigned(0 downto 0) := "0";
signal n6 : unsigned(0 downto 0) := "0";
signal n7 : unsigned(9 downto 0);
signal n8 : unsigned(9 downto 0) := "0000000000";
signal n9 : unsigned(9 downto 0) := "0000000000";
signal n10 : unsigned(9 downto 0) := "0000000000";
signal n11 : unsigned(9 downto 0) := "0000000000";
signal n12 : unsigned(0 downto 0);
signal n13 : unsigned(0 downto 0) := "0";
signal n14 : unsigned(0 downto 0) := "0";
signal n15 : unsigned(0 downto 0) := "0";
signal n16 : unsigned(0 downto 0) := "0";
signal n17 : unsigned(0 downto 0);
signal n18 : unsigned(1 downto 0);
signal n19 : unsigned(35 downto 0);
signal n20 : unsigned(35 downto 0);
signal n21 : unsigned(35 downto 0);
signal n22 : unsigned(35 downto 0);
signal n23 : unsigned(35 downto 0);
signal n24 : unsigned(35 downto 0);
signal s25_1 : unsigned(0 downto 0);
signal s26_1 : unsigned(35 downto 0);
signal s26_2 : unsigned(35 downto 0);
signal s27_1 : unsigned(10 downto 0);
signal s27_2 : unsigned(0 downto 0);
signal s28_1 : unsigned(0 downto 0);
signal s28_2 : unsigned(0 downto 0);
signal s28_3 : unsigned(71 downto 0);
signal s29_1 : unsigned(71 downto 0);
component cf_fft_4096_18_37 is
port (
clock_c : in std_logic;
i1 : in  unsigned(1 downto 0);
i2 : in  unsigned(0 downto 0);
i3 : in  unsigned(0 downto 0);
o1 : out unsigned(0 downto 0));
end component cf_fft_4096_18_37;
component cf_fft_4096_18_14 is
port (
clock_c : in std_logic;
i1 : in  unsigned(35 downto 0);
i2 : in  unsigned(35 downto 0);
i3 : in  unsigned(4 downto 0);
i4 : in  unsigned(0 downto 0);
i5 : in  unsigned(0 downto 0);
o1 : out unsigned(35 downto 0);
o2 : out unsigned(35 downto 0));
end component cf_fft_4096_18_14;
component cf_fft_4096_18_28 is
port (
clock_c : in std_logic;
i1 : in  unsigned(0 downto 0);
i2 : in  unsigned(0 downto 0);
i3 : in  unsigned(0 downto 0);
o1 : out unsigned(10 downto 0);
o2 : out unsigned(0 downto 0));
end component cf_fft_4096_18_28;
component cf_fft_4096_18_32 is
port (
clock_c : in std_logic;
i1 : in  unsigned(71 downto 0);
i2 : in  unsigned(0 downto 0);
i3 : in  unsigned(9 downto 0);
i4 : in  unsigned(0 downto 0);
i5 : in  unsigned(0 downto 0);
i6 : in  unsigned(0 downto 0);
o1 : out unsigned(0 downto 0);
o2 : out unsigned(0 downto 0);
o3 : out unsigned(71 downto 0));
end component cf_fft_4096_18_32;
component cf_fft_4096_18_33 is
port (
clock_c : in std_logic;
i1 : in  unsigned(71 downto 0);
i2 : in  unsigned(0 downto 0);
i3 : in  unsigned(9 downto 0);
i4 : in  unsigned(0 downto 0);
i5 : in  unsigned(0 downto 0);
i6 : in  unsigned(0 downto 0);
o1 : out unsigned(71 downto 0));
end component cf_fft_4096_18_33;
begin
n1 <= s27_1(10 downto 10) &
  s27_1(9 downto 9) &
  s27_1(8 downto 8) &
  s27_1(7 downto 7) &
  s27_1(6 downto 6);
n2 <= s26_1 & s26_2;
process (clock_c) begin
  if rising_edge(clock_c) then
    if i5 = "1" then
      n3 <= "0";
    elsif i4 = "1" then
      n3 <= s27_2;
    end if;
  end if;
end process;
process (clock_c) begin
  if rising_edge(clock_c) then
    if i5 = "1" then
      n4 <= "0";
    elsif i4 = "1" then
      n4 <= n3;
    end if;
  end if;
end process;
process (clock_c) begin
  if rising_edge(clock_c) then
    if i5 = "1" then
      n5 <= "0";
    elsif i4 = "1" then
      n5 <= n4;
    end if;
  end if;
end process;
process (clock_c) begin
  if rising_edge(clock_c) then
    if i5 = "1" then
      n6 <= "0";
    elsif i4 = "1" then
      n6 <= n5;
    end if;
  end if;
end process;
n7 <= s27_1(10 downto 10) &
  s27_1(9 downto 9) &
  s27_1(8 downto 8) &
  s27_1(7 downto 7) &
  s27_1(6 downto 6) &
  s27_1(5 downto 5) &
  s27_1(4 downto 4) &
  s27_1(3 downto 3) &
  s27_1(2 downto 2) &
  s27_1(1 downto 1);
process (clock_c) begin
  if rising_edge(clock_c) then
    if i5 = "1" then
      n8 <= "0000000000";
    elsif i4 = "1" then
      n8 <= n7;
    end if;
  end if;
end process;
process (clock_c) begin
  if rising_edge(clock_c) then
    if i5 = "1" then
      n9 <= "0000000000";
    elsif i4 = "1" then
      n9 <= n8;
    end if;
  end if;
end process;
process (clock_c) begin
  if rising_edge(clock_c) then
    if i5 = "1" then
      n10 <= "0000000000";
    elsif i4 = "1" then
      n10 <= n9;
    end if;
  end if;
end process;
process (clock_c) begin
  if rising_edge(clock_c) then
    if i5 = "1" then
      n11 <= "0000000000";
    elsif i4 = "1" then
      n11 <= n10;
    end if;
  end if;
end process;
n12 <= s27_1(0 downto 0);
process (clock_c) begin
  if rising_edge(clock_c) then
    if i5 = "1" then
      n13 <= "0";
    elsif i4 = "1" then
      n13 <= n12;
    end if;
  end if;
end process;
process (clock_c) begin
  if rising_edge(clock_c) then
    if i5 = "1" then
      n14 <= "0";
    elsif i4 = "1" then
      n14 <= n13;
    end if;
  end if;
end process;
process (clock_c) begin
  if rising_edge(clock_c) then
    if i5 = "1" then
      n15 <= "0";
    elsif i4 = "1" then
      n15 <= n14;
    end if;
  end if;
end process;
process (clock_c) begin
  if rising_edge(clock_c) then
    if i5 = "1" then
      n16 <= "0";
    elsif i4 = "1" then
      n16 <= n15;
    end if;
  end if;
end process;
n17 <= not n16;
n18 <= s28_2 & s28_1;
n19 <= s28_3(71 downto 71) &
  s28_3(70 downto 70) &
  s28_3(69 downto 69) &
  s28_3(68 downto 68) &
  s28_3(67 downto 67) &
  s28_3(66 downto 66) &
  s28_3(65 downto 65) &
  s28_3(64 downto 64) &
  s28_3(63 downto 63) &
  s28_3(62 downto 62) &
  s28_3(61 downto 61) &
  s28_3(60 downto 60) &
  s28_3(59 downto 59) &
  s28_3(58 downto 58) &
  s28_3(57 downto 57) &
  s28_3(56 downto 56) &
  s28_3(55 downto 55) &
  s28_3(54 downto 54) &
  s28_3(53 downto 53) &
  s28_3(52 downto 52) &
  s28_3(51 downto 51) &
  s28_3(50 downto 50) &
  s28_3(49 downto 49) &
  s28_3(48 downto 48) &
  s28_3(47 downto 47) &
  s28_3(46 downto 46) &
  s28_3(45 downto 45) &
  s28_3(44 downto 44) &
  s28_3(43 downto 43) &
  s28_3(42 downto 42) &
  s28_3(41 downto 41) &
  s28_3(40 downto 40) &
  s28_3(39 downto 39) &
  s28_3(38 downto 38) &
  s28_3(37 downto 37) &
  s28_3(36 downto 36);
n20 <= s28_3(35 downto 35) &
  s28_3(34 downto 34) &
  s28_3(33 downto 33) &
  s28_3(32 downto 32) &
  s28_3(31 downto 31) &
  s28_3(30 downto 30) &
  s28_3(29 downto 29) &
  s28_3(28 downto 28) &
  s28_3(27 downto 27) &
  s28_3(26 downto 26) &
  s28_3(25 downto 25) &
  s28_3(24 downto 24) &
  s28_3(23 downto 23) &
  s28_3(22 downto 22) &
  s28_3(21 downto 21) &
  s28_3(20 downto 20) &
  s28_3(19 downto 19) &
  s28_3(18 downto 18) &
  s28_3(17 downto 17) &
  s28_3(16 downto 16) &
  s28_3(15 downto 15) &
  s28_3(14 downto 14) &
  s28_3(13 downto 13) &
  s28_3(12 downto 12) &
  s28_3(11 downto 11) &
  s28_3(10 downto 10) &
  s28_3(9 downto 9) &
  s28_3(8 downto 8) &
  s28_3(7 downto 7) &
  s28_3(6 downto 6) &
  s28_3(5 downto 5) &
  s28_3(4 downto 4) &
  s28_3(3 downto 3) &
  s28_3(2 downto 2) &
  s28_3(1 downto 1) &
  s28_3(0 downto 0);
n21 <= s29_1(71 downto 71) &
  s29_1(70 downto 70) &
  s29_1(69 downto 69) &
  s29_1(68 downto 68) &
  s29_1(67 downto 67) &
  s29_1(66 downto 66) &
  s29_1(65 downto 65) &
  s29_1(64 downto 64) &
  s29_1(63 downto 63) &
  s29_1(62 downto 62) &
  s29_1(61 downto 61) &
  s29_1(60 downto 60) &
  s29_1(59 downto 59) &
  s29_1(58 downto 58) &
  s29_1(57 downto 57) &
  s29_1(56 downto 56) &
  s29_1(55 downto 55) &
  s29_1(54 downto 54) &
  s29_1(53 downto 53) &
  s29_1(52 downto 52) &
  s29_1(51 downto 51) &
  s29_1(50 downto 50) &
  s29_1(49 downto 49) &
  s29_1(48 downto 48) &
  s29_1(47 downto 47) &
  s29_1(46 downto 46) &
  s29_1(45 downto 45) &
  s29_1(44 downto 44) &
  s29_1(43 downto 43) &
  s29_1(42 downto 42) &
  s29_1(41 downto 41) &
  s29_1(40 downto 40) &
  s29_1(39 downto 39) &
  s29_1(38 downto 38) &
  s29_1(37 downto 37) &
  s29_1(36 downto 36);
n22 <= s29_1(35 downto 35) &
  s29_1(34 downto 34) &
  s29_1(33 downto 33) &
  s29_1(32 downto 32) &
  s29_1(31 downto 31) &
  s29_1(30 downto 30) &
  s29_1(29 downto 29) &
  s29_1(28 downto 28) &
  s29_1(27 downto 27) &
  s29_1(26 downto 26) &
  s29_1(25 downto 25) &
  s29_1(24 downto 24) &
  s29_1(23 downto 23) &
  s29_1(22 downto 22) &
  s29_1(21 downto 21) &
  s29_1(20 downto 20) &
  s29_1(19 downto 19) &
  s29_1(18 downto 18) &
  s29_1(17 downto 17) &
  s29_1(16 downto 16) &
  s29_1(15 downto 15) &
  s29_1(14 downto 14) &
  s29_1(13 downto 13) &
  s29_1(12 downto 12) &
  s29_1(11 downto 11) &
  s29_1(10 downto 10) &
  s29_1(9 downto 9) &
  s29_1(8 downto 8) &
  s29_1(7 downto 7) &
  s29_1(6 downto 6) &
  s29_1(5 downto 5) &
  s29_1(4 downto 4) &
  s29_1(3 downto 3) &
  s29_1(2 downto 2) &
  s29_1(1 downto 1) &
  s29_1(0 downto 0);
n23 <= n20 when s25_1 = "1" else n19;
n24 <= n22 when s25_1 = "1" else n21;
s25 : cf_fft_4096_18_37 port map (clock_c, n18, i4, i5, s25_1);
s26 : cf_fft_4096_18_14 port map (clock_c, i2, i3, n1, i4, i5, s26_1, s26_2);
s27 : cf_fft_4096_18_28 port map (clock_c, i1, i4, i5, s27_1, s27_2);
s28 : cf_fft_4096_18_32 port map (clock_c, n2, n6, n11, n17, i4, i5, s28_1, s28_2, s28_3);
s29 : cf_fft_4096_18_33 port map (clock_c, n2, n6, n11, n16, i4, i5, s29_1);
o3 <= n24;
o2 <= n23;
o1 <= s28_1;
end architecture rtl;

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
entity cf_fft_4096_18_12 is
port (
clock_c : in std_logic;
i1 : in  unsigned(35 downto 0);
i2 : in  unsigned(35 downto 0);
i3 : in  unsigned(3 downto 0);
i4 : in  unsigned(0 downto 0);
i5 : in  unsigned(0 downto 0);
o1 : out unsigned(35 downto 0);
o2 : out unsigned(35 downto 0));
end entity cf_fft_4096_18_12;
architecture rtl of cf_fft_4096_18_12 is
signal n1 : unsigned(35 downto 0) := "000000000000000000000000000000000000";
signal n2 : unsigned(17 downto 0);
signal n3 : unsigned(17 downto 0);
signal n4 : unsigned(35 downto 0) := "000000000000000000000000000000000000";
signal n5 : unsigned(17 downto 0);
signal n6 : unsigned(17 downto 0);
signal n7 : unsigned(17 downto 0) := "000000000000000000";
signal n8 : unsigned(17 downto 0) := "000000000000000000";
signal n9 : unsigned(17 downto 0) := "000000000000000000";
signal n10 : unsigned(17 downto 0) := "000000000000000000";
signal n11 : unsigned(35 downto 0) := "000000000000000000000000000000000000";
signal n12 : unsigned(17 downto 0);
signal n13 : unsigned(17 downto 0);
signal n14 : unsigned(35 downto 0);
signal n15 : unsigned(17 downto 0);
signal n16 : unsigned(17 downto 0) := "000000000000000000";
signal n17 : unsigned(35 downto 0);
signal n18 : unsigned(17 downto 0);
signal n19 : unsigned(17 downto 0) := "000000000000000000";
signal n20 : unsigned(17 downto 0);
signal n21 : unsigned(17 downto 0) := "000000000000000000";
signal n22 : unsigned(35 downto 0);
signal n23 : unsigned(17 downto 0);
signal n24 : unsigned(17 downto 0) := "000000000000000000";
signal n25 : unsigned(35 downto 0);
signal n26 : unsigned(17 downto 0);
signal n27 : unsigned(17 downto 0) := "000000000000000000";
signal n28 : unsigned(17 downto 0);
signal n29 : unsigned(17 downto 0) := "000000000000000000";
signal n30 : unsigned(17 downto 0);
signal n31 : unsigned(17 downto 0);
signal n32 : unsigned(35 downto 0);
signal n33 : unsigned(35 downto 0) := "000000000000000000000000000000000000";
signal n34 : unsigned(17 downto 0);
signal n35 : unsigned(17 downto 0);
signal n36 : unsigned(35 downto 0);
signal n37 : unsigned(35 downto 0) := "000000000000000000000000000000000000";
begin
process (clock_c) begin
  if rising_edge(clock_c) then
    if i5 = "1" then
      n1 <= "000000000000000000000000000000000000";
    elsif i4 = "1" then
      n1 <= i1;
    end if;
  end if;
end process;
n2 <= n1(35 downto 35) &
  n1(34 downto 34) &
  n1(33 downto 33) &
  n1(32 downto 32) &
  n1(31 downto 31) &
  n1(30 downto 30) &
  n1(29 downto 29) &
  n1(28 downto 28) &
  n1(27 downto 27) &
  n1(26 downto 26) &
  n1(25 downto 25) &
  n1(24 downto 24) &
  n1(23 downto 23) &
  n1(22 downto 22) &
  n1(21 downto 21) &
  n1(20 downto 20) &
  n1(19 downto 19) &
  n1(18 downto 18);
n3 <= n1(17 downto 17) &
  n1(16 downto 16) &
  n1(15 downto 15) &
  n1(14 downto 14) &
  n1(13 downto 13) &
  n1(12 downto 12) &
  n1(11 downto 11) &
  n1(10 downto 10) &
  n1(9 downto 9) &
  n1(8 downto 8) &
  n1(7 downto 7) &
  n1(6 downto 6) &
  n1(5 downto 5) &
  n1(4 downto 4) &
  n1(3 downto 3) &
  n1(2 downto 2) &
  n1(1 downto 1) &
  n1(0 downto 0);
process (clock_c) begin
  if rising_edge(clock_c) then
    if i5 = "1" then
      n4 <= "000000000000000000000000000000000000";
    elsif i4 = "1" then
      n4 <= i2;
    end if;
  end if;
end process;
n5 <= n4(35 downto 35) &
  n4(34 downto 34) &
  n4(33 downto 33) &
  n4(32 downto 32) &
  n4(31 downto 31) &
  n4(30 downto 30) &
  n4(29 downto 29) &
  n4(28 downto 28) &
  n4(27 downto 27) &
  n4(26 downto 26) &
  n4(25 downto 25) &
  n4(24 downto 24) &
  n4(23 downto 23) &
  n4(22 downto 22) &
  n4(21 downto 21) &
  n4(20 downto 20) &
  n4(19 downto 19) &
  n4(18 downto 18);
n6 <= n4(17 downto 17) &
  n4(16 downto 16) &
  n4(15 downto 15) &
  n4(14 downto 14) &
  n4(13 downto 13) &
  n4(12 downto 12) &
  n4(11 downto 11) &
  n4(10 downto 10) &
  n4(9 downto 9) &
  n4(8 downto 8) &
  n4(7 downto 7) &
  n4(6 downto 6) &
  n4(5 downto 5) &
  n4(4 downto 4) &
  n4(3 downto 3) &
  n4(2 downto 2) &
  n4(1 downto 1) &
  n4(0 downto 0);
process (clock_c) begin
  if rising_edge(clock_c) then
    if i5 = "1" then
      n7 <= "000000000000000000";
    elsif i4 = "1" then
      n7 <= n2;
    end if;
  end if;
end process;
process (clock_c) begin
  if rising_edge(clock_c) then
    if i5 = "1" then
      n8 <= "000000000000000000";
    elsif i4 = "1" then
      n8 <= n7;
    end if;
  end if;
end process;
process (clock_c) begin
  if rising_edge(clock_c) then
    if i5 = "1" then
      n9 <= "000000000000000000";
    elsif i4 = "1" then
      n9 <= n3;
    end if;
  end if;
end process;
process (clock_c) begin
  if rising_edge(clock_c) then
    if i5 = "1" then
      n10 <= "000000000000000000";
    elsif i4 = "1" then
      n10 <= n9;
    end if;
  end if;
end process;
process (clock_c) begin
  if rising_edge(clock_c) then 
    if i4 = "1" then
      case i3 is
        when "0000" => n11 <= "011111111111111111000000000000000000";
        when "0001" => n11 <= "011111011000101001111001110000011101";
        when "0010" => n11 <= "011101100100000110110011110000010000";
        when "0011" => n11 <= "011010100110110110101110001110001100";
        when "0100" => n11 <= "010110101000001001101001010111110110";
        when "0101" => n11 <= "010001110001110011100101011001001001";
        when "0110" => n11 <= "001100001111101111100010011011111001";
        when "0111" => n11 <= "000110001111100010100000100111010110";
        when "1000" => n11 <= "000000000000000000100000000000000000";
        when "1001" => n11 <= "111001110000011101100000100111010110";
        when "1010" => n11 <= "110011110000010000100010011011111001";
        when "1011" => n11 <= "101110001110001100100101011001001001";
        when "1100" => n11 <= "101001010111110110101001010111110110";
        when "1101" => n11 <= "100101011001001001101110001110001100";
        when "1110" => n11 <= "100010011011111001110011110000010000";
        when "1111" => n11 <= "100000100111010110111001110000011101";
        when others => n11 <= "XXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX";
      end case;
    end if;
  end if;
end process;
n12 <= n11(35 downto 35) &
  n11(34 downto 34) &
  n11(33 downto 33) &
  n11(32 downto 32) &
  n11(31 downto 31) &
  n11(30 downto 30) &
  n11(29 downto 29) &
  n11(28 downto 28) &
  n11(27 downto 27) &
  n11(26 downto 26) &
  n11(25 downto 25) &
  n11(24 downto 24) &
  n11(23 downto 23) &
  n11(22 downto 22) &
  n11(21 downto 21) &
  n11(20 downto 20) &
  n11(19 downto 19) &
  n11(18 downto 18);
n13 <= n11(17 downto 17) &
  n11(16 downto 16) &
  n11(15 downto 15) &
  n11(14 downto 14) &
  n11(13 downto 13) &
  n11(12 downto 12) &
  n11(11 downto 11) &
  n11(10 downto 10) &
  n11(9 downto 9) &
  n11(8 downto 8) &
  n11(7 downto 7) &
  n11(6 downto 6) &
  n11(5 downto 5) &
  n11(4 downto 4) &
  n11(3 downto 3) &
  n11(2 downto 2) &
  n11(1 downto 1) &
  n11(0 downto 0);
n14 <= unsigned(signed(n5) * signed(n12));
n15 <= n14(34 downto 34) &
  n14(33 downto 33) &
  n14(32 downto 32) &
  n14(31 downto 31) &
  n14(30 downto 30) &
  n14(29 downto 29) &
  n14(28 downto 28) &
  n14(27 downto 27) &
  n14(26 downto 26) &
  n14(25 downto 25) &
  n14(24 downto 24) &
  n14(23 downto 23) &
  n14(22 downto 22) &
  n14(21 downto 21) &
  n14(20 downto 20) &
  n14(19 downto 19) &
  n14(18 downto 18) &
  n14(17 downto 17);
process (clock_c) begin
  if rising_edge(clock_c) then
    if i5 = "1" then
      n16 <= "000000000000000000";
    elsif i4 = "1" then
      n16 <= n15;
    end if;
  end if;
end process;
n17 <= unsigned(signed(n6) * signed(n13));
n18 <= n17(34 downto 34) &
  n17(33 downto 33) &
  n17(32 downto 32) &
  n17(31 downto 31) &
  n17(30 downto 30) &
  n17(29 downto 29) &
  n17(28 downto 28) &
  n17(27 downto 27) &
  n17(26 downto 26) &
  n17(25 downto 25) &
  n17(24 downto 24) &
  n17(23 downto 23) &
  n17(22 downto 22) &
  n17(21 downto 21) &
  n17(20 downto 20) &
  n17(19 downto 19) &
  n17(18 downto 18) &
  n17(17 downto 17);
process (clock_c) begin
  if rising_edge(clock_c) then
    if i5 = "1" then
      n19 <= "000000000000000000";
    elsif i4 = "1" then
      n19 <= n18;
    end if;
  end if;
end process;
n20 <= n16 - n19;
process (clock_c) begin
  if rising_edge(clock_c) then
    if i5 = "1" then
      n21 <= "000000000000000000";
    elsif i4 = "1" then
      n21 <= n20;
    end if;
  end if;
end process;
n22 <= unsigned(signed(n5) * signed(n13));
n23 <= n22(34 downto 34) &
  n22(33 downto 33) &
  n22(32 downto 32) &
  n22(31 downto 31) &
  n22(30 downto 30) &
  n22(29 downto 29) &
  n22(28 downto 28) &
  n22(27 downto 27) &
  n22(26 downto 26) &
  n22(25 downto 25) &
  n22(24 downto 24) &
  n22(23 downto 23) &
  n22(22 downto 22) &
  n22(21 downto 21) &
  n22(20 downto 20) &
  n22(19 downto 19) &
  n22(18 downto 18) &
  n22(17 downto 17);
process (clock_c) begin
  if rising_edge(clock_c) then
    if i5 = "1" then
      n24 <= "000000000000000000";
    elsif i4 = "1" then
      n24 <= n23;
    end if;
  end if;
end process;
n25 <= unsigned(signed(n6) * signed(n12));
n26 <= n25(34 downto 34) &
  n25(33 downto 33) &
  n25(32 downto 32) &
  n25(31 downto 31) &
  n25(30 downto 30) &
  n25(29 downto 29) &
  n25(28 downto 28) &
  n25(27 downto 27) &
  n25(26 downto 26) &
  n25(25 downto 25) &
  n25(24 downto 24) &
  n25(23 downto 23) &
  n25(22 downto 22) &
  n25(21 downto 21) &
  n25(20 downto 20) &
  n25(19 downto 19) &
  n25(18 downto 18) &
  n25(17 downto 17);
process (clock_c) begin
  if rising_edge(clock_c) then
    if i5 = "1" then
      n27 <= "000000000000000000";
    elsif i4 = "1" then
      n27 <= n26;
    end if;
  end if;
end process;
n28 <= n24 + n27;
process (clock_c) begin
  if rising_edge(clock_c) then
    if i5 = "1" then
      n29 <= "000000000000000000";
    elsif i4 = "1" then
      n29 <= n28;
    end if;
  end if;
end process;
n30 <= n8 + n21;
n31 <= n10 + n29;
n32 <= n30 & n31;
process (clock_c) begin
  if rising_edge(clock_c) then
    if i5 = "1" then
      n33 <= "000000000000000000000000000000000000";
    elsif i4 = "1" then
      n33 <= n32;
    end if;
  end if;
end process;
n34 <= n8 - n21;
n35 <= n10 - n29;
n36 <= n34 & n35;
process (clock_c) begin
  if rising_edge(clock_c) then
    if i5 = "1" then
      n37 <= "000000000000000000000000000000000000";
    elsif i4 = "1" then
      n37 <= n36;
    end if;
  end if;
end process;
o2 <= n37;
o1 <= n33;
end architecture rtl;

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
entity cf_fft_4096_18_11 is
port (
clock_c : in std_logic;
i1 : in  unsigned(0 downto 0);
i2 : in  unsigned(35 downto 0);
i3 : in  unsigned(35 downto 0);
i4 : in  unsigned(0 downto 0);
i5 : in  unsigned(0 downto 0);
o1 : out unsigned(0 downto 0);
o2 : out unsigned(35 downto 0);
o3 : out unsigned(35 downto 0));
end entity cf_fft_4096_18_11;
architecture rtl of cf_fft_4096_18_11 is
signal n1 : unsigned(3 downto 0);
signal n2 : unsigned(71 downto 0);
signal n3 : unsigned(0 downto 0) := "0";
signal n4 : unsigned(0 downto 0) := "0";
signal n5 : unsigned(0 downto 0) := "0";
signal n6 : unsigned(0 downto 0) := "0";
signal n7 : unsigned(9 downto 0);
signal n8 : unsigned(9 downto 0) := "0000000000";
signal n9 : unsigned(9 downto 0) := "0000000000";
signal n10 : unsigned(9 downto 0) := "0000000000";
signal n11 : unsigned(9 downto 0) := "0000000000";
signal n12 : unsigned(0 downto 0);
signal n13 : unsigned(0 downto 0) := "0";
signal n14 : unsigned(0 downto 0) := "0";
signal n15 : unsigned(0 downto 0) := "0";
signal n16 : unsigned(0 downto 0) := "0";
signal n17 : unsigned(0 downto 0);
signal n18 : unsigned(1 downto 0);
signal n19 : unsigned(35 downto 0);
signal n20 : unsigned(35 downto 0);
signal n21 : unsigned(35 downto 0);
signal n22 : unsigned(35 downto 0);
signal n23 : unsigned(35 downto 0);
signal n24 : unsigned(35 downto 0);
signal s25_1 : unsigned(35 downto 0);
signal s25_2 : unsigned(35 downto 0);
signal s26_1 : unsigned(0 downto 0);
signal s27_1 : unsigned(0 downto 0);
signal s27_2 : unsigned(0 downto 0);
signal s27_3 : unsigned(71 downto 0);
signal s28_1 : unsigned(71 downto 0);
signal s29_1 : unsigned(10 downto 0);
signal s29_2 : unsigned(0 downto 0);
component cf_fft_4096_18_12 is
port (
clock_c : in std_logic;
i1 : in  unsigned(35 downto 0);
i2 : in  unsigned(35 downto 0);
i3 : in  unsigned(3 downto 0);
i4 : in  unsigned(0 downto 0);
i5 : in  unsigned(0 downto 0);
o1 : out unsigned(35 downto 0);
o2 : out unsigned(35 downto 0));
end component cf_fft_4096_18_12;
component cf_fft_4096_18_37 is
port (
clock_c : in std_logic;
i1 : in  unsigned(1 downto 0);
i2 : in  unsigned(0 downto 0);
i3 : in  unsigned(0 downto 0);
o1 : out unsigned(0 downto 0));
end component cf_fft_4096_18_37;
component cf_fft_4096_18_32 is
port (
clock_c : in std_logic;
i1 : in  unsigned(71 downto 0);
i2 : in  unsigned(0 downto 0);
i3 : in  unsigned(9 downto 0);
i4 : in  unsigned(0 downto 0);
i5 : in  unsigned(0 downto 0);
i6 : in  unsigned(0 downto 0);
o1 : out unsigned(0 downto 0);
o2 : out unsigned(0 downto 0);
o3 : out unsigned(71 downto 0));
end component cf_fft_4096_18_32;
component cf_fft_4096_18_33 is
port (
clock_c : in std_logic;
i1 : in  unsigned(71 downto 0);
i2 : in  unsigned(0 downto 0);
i3 : in  unsigned(9 downto 0);
i4 : in  unsigned(0 downto 0);
i5 : in  unsigned(0 downto 0);
i6 : in  unsigned(0 downto 0);
o1 : out unsigned(71 downto 0));
end component cf_fft_4096_18_33;
component cf_fft_4096_18_28 is
port (
clock_c : in std_logic;
i1 : in  unsigned(0 downto 0);
i2 : in  unsigned(0 downto 0);
i3 : in  unsigned(0 downto 0);
o1 : out unsigned(10 downto 0);
o2 : out unsigned(0 downto 0));
end component cf_fft_4096_18_28;
begin
n1 <= s29_1(10 downto 10) &
  s29_1(9 downto 9) &
  s29_1(8 downto 8) &
  s29_1(7 downto 7);
n2 <= s25_1 & s25_2;
process (clock_c) begin
  if rising_edge(clock_c) then
    if i5 = "1" then
      n3 <= "0";
    elsif i4 = "1" then
      n3 <= s29_2;
    end if;
  end if;
end process;
process (clock_c) begin
  if rising_edge(clock_c) then
    if i5 = "1" then
      n4 <= "0";
    elsif i4 = "1" then
      n4 <= n3;
    end if;
  end if;
end process;
process (clock_c) begin
  if rising_edge(clock_c) then
    if i5 = "1" then
      n5 <= "0";
    elsif i4 = "1" then
      n5 <= n4;
    end if;
  end if;
end process;
process (clock_c) begin
  if rising_edge(clock_c) then
    if i5 = "1" then
      n6 <= "0";
    elsif i4 = "1" then
      n6 <= n5;
    end if;
  end if;
end process;
n7 <= s29_1(10 downto 10) &
  s29_1(9 downto 9) &
  s29_1(8 downto 8) &
  s29_1(7 downto 7) &
  s29_1(6 downto 6) &
  s29_1(5 downto 5) &
  s29_1(4 downto 4) &
  s29_1(3 downto 3) &
  s29_1(2 downto 2) &
  s29_1(1 downto 1);
process (clock_c) begin
  if rising_edge(clock_c) then
    if i5 = "1" then
      n8 <= "0000000000";
    elsif i4 = "1" then
      n8 <= n7;
    end if;
  end if;
end process;
process (clock_c) begin
  if rising_edge(clock_c) then
    if i5 = "1" then
      n9 <= "0000000000";
    elsif i4 = "1" then
      n9 <= n8;
    end if;
  end if;
end process;
process (clock_c) begin
  if rising_edge(clock_c) then
    if i5 = "1" then
      n10 <= "0000000000";
    elsif i4 = "1" then
      n10 <= n9;
    end if;
  end if;
end process;
process (clock_c) begin
  if rising_edge(clock_c) then
    if i5 = "1" then
      n11 <= "0000000000";
    elsif i4 = "1" then
      n11 <= n10;
    end if;
  end if;
end process;
n12 <= s29_1(0 downto 0);
process (clock_c) begin
  if rising_edge(clock_c) then
    if i5 = "1" then
      n13 <= "0";
    elsif i4 = "1" then
      n13 <= n12;
    end if;
  end if;
end process;
process (clock_c) begin
  if rising_edge(clock_c) then
    if i5 = "1" then
      n14 <= "0";
    elsif i4 = "1" then
      n14 <= n13;
    end if;
  end if;
end process;
process (clock_c) begin
  if rising_edge(clock_c) then
    if i5 = "1" then
      n15 <= "0";
    elsif i4 = "1" then
      n15 <= n14;
    end if;
  end if;
end process;
process (clock_c) begin
  if rising_edge(clock_c) then
    if i5 = "1" then
      n16 <= "0";
    elsif i4 = "1" then
      n16 <= n15;
    end if;
  end if;
end process;
n17 <= not n16;
n18 <= s27_2 & s27_1;
n19 <= s27_3(71 downto 71) &
  s27_3(70 downto 70) &
  s27_3(69 downto 69) &
  s27_3(68 downto 68) &
  s27_3(67 downto 67) &
  s27_3(66 downto 66) &
  s27_3(65 downto 65) &
  s27_3(64 downto 64) &
  s27_3(63 downto 63) &
  s27_3(62 downto 62) &
  s27_3(61 downto 61) &
  s27_3(60 downto 60) &
  s27_3(59 downto 59) &
  s27_3(58 downto 58) &
  s27_3(57 downto 57) &
  s27_3(56 downto 56) &
  s27_3(55 downto 55) &
  s27_3(54 downto 54) &
  s27_3(53 downto 53) &
  s27_3(52 downto 52) &
  s27_3(51 downto 51) &
  s27_3(50 downto 50) &
  s27_3(49 downto 49) &
  s27_3(48 downto 48) &
  s27_3(47 downto 47) &
  s27_3(46 downto 46) &
  s27_3(45 downto 45) &
  s27_3(44 downto 44) &
  s27_3(43 downto 43) &
  s27_3(42 downto 42) &
  s27_3(41 downto 41) &
  s27_3(40 downto 40) &
  s27_3(39 downto 39) &
  s27_3(38 downto 38) &
  s27_3(37 downto 37) &
  s27_3(36 downto 36);
n20 <= s27_3(35 downto 35) &
  s27_3(34 downto 34) &
  s27_3(33 downto 33) &
  s27_3(32 downto 32) &
  s27_3(31 downto 31) &
  s27_3(30 downto 30) &
  s27_3(29 downto 29) &
  s27_3(28 downto 28) &
  s27_3(27 downto 27) &
  s27_3(26 downto 26) &
  s27_3(25 downto 25) &
  s27_3(24 downto 24) &
  s27_3(23 downto 23) &
  s27_3(22 downto 22) &
  s27_3(21 downto 21) &
  s27_3(20 downto 20) &
  s27_3(19 downto 19) &
  s27_3(18 downto 18) &
  s27_3(17 downto 17) &
  s27_3(16 downto 16) &
  s27_3(15 downto 15) &
  s27_3(14 downto 14) &
  s27_3(13 downto 13) &
  s27_3(12 downto 12) &
  s27_3(11 downto 11) &
  s27_3(10 downto 10) &
  s27_3(9 downto 9) &
  s27_3(8 downto 8) &
  s27_3(7 downto 7) &
  s27_3(6 downto 6) &
  s27_3(5 downto 5) &
  s27_3(4 downto 4) &
  s27_3(3 downto 3) &
  s27_3(2 downto 2) &
  s27_3(1 downto 1) &
  s27_3(0 downto 0);
n21 <= s28_1(71 downto 71) &
  s28_1(70 downto 70) &
  s28_1(69 downto 69) &
  s28_1(68 downto 68) &
  s28_1(67 downto 67) &
  s28_1(66 downto 66) &
  s28_1(65 downto 65) &
  s28_1(64 downto 64) &
  s28_1(63 downto 63) &
  s28_1(62 downto 62) &
  s28_1(61 downto 61) &
  s28_1(60 downto 60) &
  s28_1(59 downto 59) &
  s28_1(58 downto 58) &
  s28_1(57 downto 57) &
  s28_1(56 downto 56) &
  s28_1(55 downto 55) &
  s28_1(54 downto 54) &
  s28_1(53 downto 53) &
  s28_1(52 downto 52) &
  s28_1(51 downto 51) &
  s28_1(50 downto 50) &
  s28_1(49 downto 49) &
  s28_1(48 downto 48) &
  s28_1(47 downto 47) &
  s28_1(46 downto 46) &
  s28_1(45 downto 45) &
  s28_1(44 downto 44) &
  s28_1(43 downto 43) &
  s28_1(42 downto 42) &
  s28_1(41 downto 41) &
  s28_1(40 downto 40) &
  s28_1(39 downto 39) &
  s28_1(38 downto 38) &
  s28_1(37 downto 37) &
  s28_1(36 downto 36);
n22 <= s28_1(35 downto 35) &
  s28_1(34 downto 34) &
  s28_1(33 downto 33) &
  s28_1(32 downto 32) &
  s28_1(31 downto 31) &
  s28_1(30 downto 30) &
  s28_1(29 downto 29) &
  s28_1(28 downto 28) &
  s28_1(27 downto 27) &
  s28_1(26 downto 26) &
  s28_1(25 downto 25) &
  s28_1(24 downto 24) &
  s28_1(23 downto 23) &
  s28_1(22 downto 22) &
  s28_1(21 downto 21) &
  s28_1(20 downto 20) &
  s28_1(19 downto 19) &
  s28_1(18 downto 18) &
  s28_1(17 downto 17) &
  s28_1(16 downto 16) &
  s28_1(15 downto 15) &
  s28_1(14 downto 14) &
  s28_1(13 downto 13) &
  s28_1(12 downto 12) &
  s28_1(11 downto 11) &
  s28_1(10 downto 10) &
  s28_1(9 downto 9) &
  s28_1(8 downto 8) &
  s28_1(7 downto 7) &
  s28_1(6 downto 6) &
  s28_1(5 downto 5) &
  s28_1(4 downto 4) &
  s28_1(3 downto 3) &
  s28_1(2 downto 2) &
  s28_1(1 downto 1) &
  s28_1(0 downto 0);
n23 <= n20 when s26_1 = "1" else n19;
n24 <= n22 when s26_1 = "1" else n21;
s25 : cf_fft_4096_18_12 port map (clock_c, i2, i3, n1, i4, i5, s25_1, s25_2);
s26 : cf_fft_4096_18_37 port map (clock_c, n18, i4, i5, s26_1);
s27 : cf_fft_4096_18_32 port map (clock_c, n2, n6, n11, n17, i4, i5, s27_1, s27_2, s27_3);
s28 : cf_fft_4096_18_33 port map (clock_c, n2, n6, n11, n16, i4, i5, s28_1);
s29 : cf_fft_4096_18_28 port map (clock_c, i1, i4, i5, s29_1, s29_2);
o3 <= n24;
o2 <= n23;
o1 <= s27_1;
end architecture rtl;

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
entity cf_fft_4096_18_10 is
port (
clock_c : in std_logic;
i1 : in  unsigned(0 downto 0);
i2 : in  unsigned(35 downto 0);
i3 : in  unsigned(35 downto 0);
i4 : in  unsigned(0 downto 0);
i5 : in  unsigned(0 downto 0);
o1 : out unsigned(0 downto 0);
o2 : out unsigned(35 downto 0);
o3 : out unsigned(35 downto 0));
end entity cf_fft_4096_18_10;
architecture rtl of cf_fft_4096_18_10 is
signal s1_1 : unsigned(0 downto 0);
signal s1_2 : unsigned(35 downto 0);
signal s1_3 : unsigned(35 downto 0);
signal s2_1 : unsigned(0 downto 0);
signal s2_2 : unsigned(35 downto 0);
signal s2_3 : unsigned(35 downto 0);
signal s3_1 : unsigned(0 downto 0);
signal s3_2 : unsigned(35 downto 0);
signal s3_3 : unsigned(35 downto 0);
signal s4_1 : unsigned(0 downto 0);
signal s4_2 : unsigned(35 downto 0);
signal s4_3 : unsigned(35 downto 0);
signal s5_1 : unsigned(0 downto 0);
signal s5_2 : unsigned(35 downto 0);
signal s5_3 : unsigned(35 downto 0);
signal s6_1 : unsigned(0 downto 0);
signal s6_2 : unsigned(35 downto 0);
signal s6_3 : unsigned(35 downto 0);
signal s7_1 : unsigned(0 downto 0);
signal s7_2 : unsigned(35 downto 0);
signal s7_3 : unsigned(35 downto 0);
signal s8_1 : unsigned(0 downto 0);
signal s8_2 : unsigned(35 downto 0);
signal s8_3 : unsigned(35 downto 0);
component cf_fft_4096_18_25 is
port (
clock_c : in std_logic;
i1 : in  unsigned(0 downto 0);
i2 : in  unsigned(35 downto 0);
i3 : in  unsigned(35 downto 0);
i4 : in  unsigned(0 downto 0);
i5 : in  unsigned(0 downto 0);
o1 : out unsigned(0 downto 0);
o2 : out unsigned(35 downto 0);
o3 : out unsigned(35 downto 0));
end component cf_fft_4096_18_25;
component cf_fft_4096_18_23 is
port (
clock_c : in std_logic;
i1 : in  unsigned(0 downto 0);
i2 : in  unsigned(35 downto 0);
i3 : in  unsigned(35 downto 0);
i4 : in  unsigned(0 downto 0);
i5 : in  unsigned(0 downto 0);
o1 : out unsigned(0 downto 0);
o2 : out unsigned(35 downto 0);
o3 : out unsigned(35 downto 0));
end component cf_fft_4096_18_23;
component cf_fft_4096_18_21 is
port (
clock_c : in std_logic;
i1 : in  unsigned(0 downto 0);
i2 : in  unsigned(35 downto 0);
i3 : in  unsigned(35 downto 0);
i4 : in  unsigned(0 downto 0);
i5 : in  unsigned(0 downto 0);
o1 : out unsigned(0 downto 0);
o2 : out unsigned(35 downto 0);
o3 : out unsigned(35 downto 0));
end component cf_fft_4096_18_21;
component cf_fft_4096_18_19 is
port (
clock_c : in std_logic;
i1 : in  unsigned(0 downto 0);
i2 : in  unsigned(35 downto 0);
i3 : in  unsigned(35 downto 0);
i4 : in  unsigned(0 downto 0);
i5 : in  unsigned(0 downto 0);
o1 : out unsigned(0 downto 0);
o2 : out unsigned(35 downto 0);
o3 : out unsigned(35 downto 0));
end component cf_fft_4096_18_19;
component cf_fft_4096_18_17 is
port (
clock_c : in std_logic;
i1 : in  unsigned(0 downto 0);
i2 : in  unsigned(35 downto 0);
i3 : in  unsigned(35 downto 0);
i4 : in  unsigned(0 downto 0);
i5 : in  unsigned(0 downto 0);
o1 : out unsigned(0 downto 0);
o2 : out unsigned(35 downto 0);
o3 : out unsigned(35 downto 0));
end component cf_fft_4096_18_17;
component cf_fft_4096_18_15 is
port (
clock_c : in std_logic;
i1 : in  unsigned(0 downto 0);
i2 : in  unsigned(35 downto 0);
i3 : in  unsigned(35 downto 0);
i4 : in  unsigned(0 downto 0);
i5 : in  unsigned(0 downto 0);
o1 : out unsigned(0 downto 0);
o2 : out unsigned(35 downto 0);
o3 : out unsigned(35 downto 0));
end component cf_fft_4096_18_15;
component cf_fft_4096_18_13 is
port (
clock_c : in std_logic;
i1 : in  unsigned(0 downto 0);
i2 : in  unsigned(35 downto 0);
i3 : in  unsigned(35 downto 0);
i4 : in  unsigned(0 downto 0);
i5 : in  unsigned(0 downto 0);
o1 : out unsigned(0 downto 0);
o2 : out unsigned(35 downto 0);
o3 : out unsigned(35 downto 0));
end component cf_fft_4096_18_13;
component cf_fft_4096_18_11 is
port (
clock_c : in std_logic;
i1 : in  unsigned(0 downto 0);
i2 : in  unsigned(35 downto 0);
i3 : in  unsigned(35 downto 0);
i4 : in  unsigned(0 downto 0);
i5 : in  unsigned(0 downto 0);
o1 : out unsigned(0 downto 0);
o2 : out unsigned(35 downto 0);
o3 : out unsigned(35 downto 0));
end component cf_fft_4096_18_11;
begin
s1 : cf_fft_4096_18_25 port map (clock_c, s2_1, s2_2, s2_3, i4, i5, s1_1, s1_2, s1_3);
s2 : cf_fft_4096_18_23 port map (clock_c, s3_1, s3_2, s3_3, i4, i5, s2_1, s2_2, s2_3);
s3 : cf_fft_4096_18_21 port map (clock_c, s4_1, s4_2, s4_3, i4, i5, s3_1, s3_2, s3_3);
s4 : cf_fft_4096_18_19 port map (clock_c, s5_1, s5_2, s5_3, i4, i5, s4_1, s4_2, s4_3);
s5 : cf_fft_4096_18_17 port map (clock_c, s6_1, s6_2, s6_3, i4, i5, s5_1, s5_2, s5_3);
s6 : cf_fft_4096_18_15 port map (clock_c, s7_1, s7_2, s7_3, i4, i5, s6_1, s6_2, s6_3);
s7 : cf_fft_4096_18_13 port map (clock_c, s8_1, s8_2, s8_3, i4, i5, s7_1, s7_2, s7_3);
s8 : cf_fft_4096_18_11 port map (clock_c, i1, i2, i3, i4, i5, s8_1, s8_2, s8_3);
o3 <= s1_3;
o2 <= s1_2;
o1 <= s1_1;
end architecture rtl;

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
entity cf_fft_4096_18_9 is
port (
clock_c : in std_logic;
i1 : in  unsigned(35 downto 0);
i2 : in  unsigned(35 downto 0);
i3 : in  unsigned(1 downto 0);
i4 : in  unsigned(0 downto 0);
i5 : in  unsigned(0 downto 0);
o1 : out unsigned(35 downto 0);
o2 : out unsigned(35 downto 0));
end entity cf_fft_4096_18_9;
architecture rtl of cf_fft_4096_18_9 is
signal n1 : unsigned(35 downto 0) := "000000000000000000000000000000000000";
signal n2 : unsigned(17 downto 0);
signal n3 : unsigned(17 downto 0);
signal n4 : unsigned(35 downto 0) := "000000000000000000000000000000000000";
signal n5 : unsigned(17 downto 0);
signal n6 : unsigned(17 downto 0);
signal n7 : unsigned(17 downto 0) := "000000000000000000";
signal n8 : unsigned(17 downto 0) := "000000000000000000";
signal n9 : unsigned(17 downto 0) := "000000000000000000";
signal n10 : unsigned(17 downto 0) := "000000000000000000";
signal n11 : unsigned(35 downto 0) := "000000000000000000000000000000000000";
signal n12 : unsigned(17 downto 0);
signal n13 : unsigned(17 downto 0);
signal n14 : unsigned(35 downto 0);
signal n15 : unsigned(17 downto 0);
signal n16 : unsigned(17 downto 0) := "000000000000000000";
signal n17 : unsigned(35 downto 0);
signal n18 : unsigned(17 downto 0);
signal n19 : unsigned(17 downto 0) := "000000000000000000";
signal n20 : unsigned(17 downto 0);
signal n21 : unsigned(17 downto 0) := "000000000000000000";
signal n22 : unsigned(35 downto 0);
signal n23 : unsigned(17 downto 0);
signal n24 : unsigned(17 downto 0) := "000000000000000000";
signal n25 : unsigned(35 downto 0);
signal n26 : unsigned(17 downto 0);
signal n27 : unsigned(17 downto 0) := "000000000000000000";
signal n28 : unsigned(17 downto 0);
signal n29 : unsigned(17 downto 0) := "000000000000000000";
signal n30 : unsigned(17 downto 0);
signal n31 : unsigned(17 downto 0);
signal n32 : unsigned(35 downto 0);
signal n33 : unsigned(35 downto 0) := "000000000000000000000000000000000000";
signal n34 : unsigned(17 downto 0);
signal n35 : unsigned(17 downto 0);
signal n36 : unsigned(35 downto 0);
signal n37 : unsigned(35 downto 0) := "000000000000000000000000000000000000";
begin
process (clock_c) begin
  if rising_edge(clock_c) then
    if i5 = "1" then
      n1 <= "000000000000000000000000000000000000";
    elsif i4 = "1" then
      n1 <= i1;
    end if;
  end if;
end process;
n2 <= n1(35 downto 35) &
  n1(34 downto 34) &
  n1(33 downto 33) &
  n1(32 downto 32) &
  n1(31 downto 31) &
  n1(30 downto 30) &
  n1(29 downto 29) &
  n1(28 downto 28) &
  n1(27 downto 27) &
  n1(26 downto 26) &
  n1(25 downto 25) &
  n1(24 downto 24) &
  n1(23 downto 23) &
  n1(22 downto 22) &
  n1(21 downto 21) &
  n1(20 downto 20) &
  n1(19 downto 19) &
  n1(18 downto 18);
n3 <= n1(17 downto 17) &
  n1(16 downto 16) &
  n1(15 downto 15) &
  n1(14 downto 14) &
  n1(13 downto 13) &
  n1(12 downto 12) &
  n1(11 downto 11) &
  n1(10 downto 10) &
  n1(9 downto 9) &
  n1(8 downto 8) &
  n1(7 downto 7) &
  n1(6 downto 6) &
  n1(5 downto 5) &
  n1(4 downto 4) &
  n1(3 downto 3) &
  n1(2 downto 2) &
  n1(1 downto 1) &
  n1(0 downto 0);
process (clock_c) begin
  if rising_edge(clock_c) then
    if i5 = "1" then
      n4 <= "000000000000000000000000000000000000";
    elsif i4 = "1" then
      n4 <= i2;
    end if;
  end if;
end process;
n5 <= n4(35 downto 35) &
  n4(34 downto 34) &
  n4(33 downto 33) &
  n4(32 downto 32) &
  n4(31 downto 31) &
  n4(30 downto 30) &
  n4(29 downto 29) &
  n4(28 downto 28) &
  n4(27 downto 27) &
  n4(26 downto 26) &
  n4(25 downto 25) &
  n4(24 downto 24) &
  n4(23 downto 23) &
  n4(22 downto 22) &
  n4(21 downto 21) &
  n4(20 downto 20) &
  n4(19 downto 19) &
  n4(18 downto 18);
n6 <= n4(17 downto 17) &
  n4(16 downto 16) &
  n4(15 downto 15) &
  n4(14 downto 14) &
  n4(13 downto 13) &
  n4(12 downto 12) &
  n4(11 downto 11) &
  n4(10 downto 10) &
  n4(9 downto 9) &
  n4(8 downto 8) &
  n4(7 downto 7) &
  n4(6 downto 6) &
  n4(5 downto 5) &
  n4(4 downto 4) &
  n4(3 downto 3) &
  n4(2 downto 2) &
  n4(1 downto 1) &
  n4(0 downto 0);
process (clock_c) begin
  if rising_edge(clock_c) then
    if i5 = "1" then
      n7 <= "000000000000000000";
    elsif i4 = "1" then
      n7 <= n2;
    end if;
  end if;
end process;
process (clock_c) begin
  if rising_edge(clock_c) then
    if i5 = "1" then
      n8 <= "000000000000000000";
    elsif i4 = "1" then
      n8 <= n7;
    end if;
  end if;
end process;
process (clock_c) begin
  if rising_edge(clock_c) then
    if i5 = "1" then
      n9 <= "000000000000000000";
    elsif i4 = "1" then
      n9 <= n3;
    end if;
  end if;
end process;
process (clock_c) begin
  if rising_edge(clock_c) then
    if i5 = "1" then
      n10 <= "000000000000000000";
    elsif i4 = "1" then
      n10 <= n9;
    end if;
  end if;
end process;
process (clock_c) begin
  if rising_edge(clock_c) then 
    if i4 = "1" then
      case i3 is
        when "00" => n11 <= "011111111111111111000000000000000000";
        when "01" => n11 <= "010110101000001001101001010111110110";
        when "10" => n11 <= "000000000000000000100000000000000000";
        when "11" => n11 <= "101001010111110110101001010111110110";
        when others => n11 <= "XXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX";
      end case;
    end if;
  end if;
end process;
n12 <= n11(35 downto 35) &
  n11(34 downto 34) &
  n11(33 downto 33) &
  n11(32 downto 32) &
  n11(31 downto 31) &
  n11(30 downto 30) &
  n11(29 downto 29) &
  n11(28 downto 28) &
  n11(27 downto 27) &
  n11(26 downto 26) &
  n11(25 downto 25) &
  n11(24 downto 24) &
  n11(23 downto 23) &
  n11(22 downto 22) &
  n11(21 downto 21) &
  n11(20 downto 20) &
  n11(19 downto 19) &
  n11(18 downto 18);
n13 <= n11(17 downto 17) &
  n11(16 downto 16) &
  n11(15 downto 15) &
  n11(14 downto 14) &
  n11(13 downto 13) &
  n11(12 downto 12) &
  n11(11 downto 11) &
  n11(10 downto 10) &
  n11(9 downto 9) &
  n11(8 downto 8) &
  n11(7 downto 7) &
  n11(6 downto 6) &
  n11(5 downto 5) &
  n11(4 downto 4) &
  n11(3 downto 3) &
  n11(2 downto 2) &
  n11(1 downto 1) &
  n11(0 downto 0);
n14 <= unsigned(signed(n5) * signed(n12));
n15 <= n14(34 downto 34) &
  n14(33 downto 33) &
  n14(32 downto 32) &
  n14(31 downto 31) &
  n14(30 downto 30) &
  n14(29 downto 29) &
  n14(28 downto 28) &
  n14(27 downto 27) &
  n14(26 downto 26) &
  n14(25 downto 25) &
  n14(24 downto 24) &
  n14(23 downto 23) &
  n14(22 downto 22) &
  n14(21 downto 21) &
  n14(20 downto 20) &
  n14(19 downto 19) &
  n14(18 downto 18) &
  n14(17 downto 17);
process (clock_c) begin
  if rising_edge(clock_c) then
    if i5 = "1" then
      n16 <= "000000000000000000";
    elsif i4 = "1" then
      n16 <= n15;
    end if;
  end if;
end process;
n17 <= unsigned(signed(n6) * signed(n13));
n18 <= n17(34 downto 34) &
  n17(33 downto 33) &
  n17(32 downto 32) &
  n17(31 downto 31) &
  n17(30 downto 30) &
  n17(29 downto 29) &
  n17(28 downto 28) &
  n17(27 downto 27) &
  n17(26 downto 26) &
  n17(25 downto 25) &
  n17(24 downto 24) &
  n17(23 downto 23) &
  n17(22 downto 22) &
  n17(21 downto 21) &
  n17(20 downto 20) &
  n17(19 downto 19) &
  n17(18 downto 18) &
  n17(17 downto 17);
process (clock_c) begin
  if rising_edge(clock_c) then
    if i5 = "1" then
      n19 <= "000000000000000000";
    elsif i4 = "1" then
      n19 <= n18;
    end if;
  end if;
end process;
n20 <= n16 - n19;
process (clock_c) begin
  if rising_edge(clock_c) then
    if i5 = "1" then
      n21 <= "000000000000000000";
    elsif i4 = "1" then
      n21 <= n20;
    end if;
  end if;
end process;
n22 <= unsigned(signed(n5) * signed(n13));
n23 <= n22(34 downto 34) &
  n22(33 downto 33) &
  n22(32 downto 32) &
  n22(31 downto 31) &
  n22(30 downto 30) &
  n22(29 downto 29) &
  n22(28 downto 28) &
  n22(27 downto 27) &
  n22(26 downto 26) &
  n22(25 downto 25) &
  n22(24 downto 24) &
  n22(23 downto 23) &
  n22(22 downto 22) &
  n22(21 downto 21) &
  n22(20 downto 20) &
  n22(19 downto 19) &
  n22(18 downto 18) &
  n22(17 downto 17);
process (clock_c) begin
  if rising_edge(clock_c) then
    if i5 = "1" then
      n24 <= "000000000000000000";
    elsif i4 = "1" then
      n24 <= n23;
    end if;
  end if;
end process;
n25 <= unsigned(signed(n6) * signed(n12));
n26 <= n25(34 downto 34) &
  n25(33 downto 33) &
  n25(32 downto 32) &
  n25(31 downto 31) &
  n25(30 downto 30) &
  n25(29 downto 29) &
  n25(28 downto 28) &
  n25(27 downto 27) &
  n25(26 downto 26) &
  n25(25 downto 25) &
  n25(24 downto 24) &
  n25(23 downto 23) &
  n25(22 downto 22) &
  n25(21 downto 21) &
  n25(20 downto 20) &
  n25(19 downto 19) &
  n25(18 downto 18) &
  n25(17 downto 17);
process (clock_c) begin
  if rising_edge(clock_c) then
    if i5 = "1" then
      n27 <= "000000000000000000";
    elsif i4 = "1" then
      n27 <= n26;
    end if;
  end if;
end process;
n28 <= n24 + n27;
process (clock_c) begin
  if rising_edge(clock_c) then
    if i5 = "1" then
      n29 <= "000000000000000000";
    elsif i4 = "1" then
      n29 <= n28;
    end if;
  end if;
end process;
n30 <= n8 + n21;
n31 <= n10 + n29;
n32 <= n30 & n31;
process (clock_c) begin
  if rising_edge(clock_c) then
    if i5 = "1" then
      n33 <= "000000000000000000000000000000000000";
    elsif i4 = "1" then
      n33 <= n32;
    end if;
  end if;
end process;
n34 <= n8 - n21;
n35 <= n10 - n29;
n36 <= n34 & n35;
process (clock_c) begin
  if rising_edge(clock_c) then
    if i5 = "1" then
      n37 <= "000000000000000000000000000000000000";
    elsif i4 = "1" then
      n37 <= n36;
    end if;
  end if;
end process;
o2 <= n37;
o1 <= n33;
end architecture rtl;

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
entity cf_fft_4096_18_8 is
port (
clock_c : in std_logic;
i1 : in  unsigned(0 downto 0);
i2 : in  unsigned(35 downto 0);
i3 : in  unsigned(35 downto 0);
i4 : in  unsigned(0 downto 0);
i5 : in  unsigned(0 downto 0);
o1 : out unsigned(0 downto 0);
o2 : out unsigned(35 downto 0);
o3 : out unsigned(35 downto 0));
end entity cf_fft_4096_18_8;
architecture rtl of cf_fft_4096_18_8 is
signal n1 : unsigned(1 downto 0);
signal n2 : unsigned(71 downto 0);
signal n3 : unsigned(0 downto 0) := "0";
signal n4 : unsigned(0 downto 0) := "0";
signal n5 : unsigned(0 downto 0) := "0";
signal n6 : unsigned(0 downto 0) := "0";
signal n7 : unsigned(9 downto 0);
signal n8 : unsigned(9 downto 0) := "0000000000";
signal n9 : unsigned(9 downto 0) := "0000000000";
signal n10 : unsigned(9 downto 0) := "0000000000";
signal n11 : unsigned(9 downto 0) := "0000000000";
signal n12 : unsigned(0 downto 0);
signal n13 : unsigned(0 downto 0) := "0";
signal n14 : unsigned(0 downto 0) := "0";
signal n15 : unsigned(0 downto 0) := "0";
signal n16 : unsigned(0 downto 0) := "0";
signal n17 : unsigned(0 downto 0);
signal n18 : unsigned(1 downto 0);
signal n19 : unsigned(35 downto 0);
signal n20 : unsigned(35 downto 0);
signal n21 : unsigned(35 downto 0);
signal n22 : unsigned(35 downto 0);
signal n23 : unsigned(35 downto 0);
signal n24 : unsigned(35 downto 0);
signal s25_1 : unsigned(35 downto 0);
signal s25_2 : unsigned(35 downto 0);
signal s26_1 : unsigned(0 downto 0);
signal s27_1 : unsigned(71 downto 0);
signal s28_1 : unsigned(0 downto 0);
signal s28_2 : unsigned(0 downto 0);
signal s28_3 : unsigned(71 downto 0);
signal s29_1 : unsigned(10 downto 0);
signal s29_2 : unsigned(0 downto 0);
component cf_fft_4096_18_9 is
port (
clock_c : in std_logic;
i1 : in  unsigned(35 downto 0);
i2 : in  unsigned(35 downto 0);
i3 : in  unsigned(1 downto 0);
i4 : in  unsigned(0 downto 0);
i5 : in  unsigned(0 downto 0);
o1 : out unsigned(35 downto 0);
o2 : out unsigned(35 downto 0));
end component cf_fft_4096_18_9;
component cf_fft_4096_18_37 is
port (
clock_c : in std_logic;
i1 : in  unsigned(1 downto 0);
i2 : in  unsigned(0 downto 0);
i3 : in  unsigned(0 downto 0);
o1 : out unsigned(0 downto 0));
end component cf_fft_4096_18_37;
component cf_fft_4096_18_33 is
port (
clock_c : in std_logic;
i1 : in  unsigned(71 downto 0);
i2 : in  unsigned(0 downto 0);
i3 : in  unsigned(9 downto 0);
i4 : in  unsigned(0 downto 0);
i5 : in  unsigned(0 downto 0);
i6 : in  unsigned(0 downto 0);
o1 : out unsigned(71 downto 0));
end component cf_fft_4096_18_33;
component cf_fft_4096_18_32 is
port (
clock_c : in std_logic;
i1 : in  unsigned(71 downto 0);
i2 : in  unsigned(0 downto 0);
i3 : in  unsigned(9 downto 0);
i4 : in  unsigned(0 downto 0);
i5 : in  unsigned(0 downto 0);
i6 : in  unsigned(0 downto 0);
o1 : out unsigned(0 downto 0);
o2 : out unsigned(0 downto 0);
o3 : out unsigned(71 downto 0));
end component cf_fft_4096_18_32;
component cf_fft_4096_18_28 is
port (
clock_c : in std_logic;
i1 : in  unsigned(0 downto 0);
i2 : in  unsigned(0 downto 0);
i3 : in  unsigned(0 downto 0);
o1 : out unsigned(10 downto 0);
o2 : out unsigned(0 downto 0));
end component cf_fft_4096_18_28;
begin
n1 <= s29_1(10 downto 10) &
  s29_1(9 downto 9);
n2 <= s25_1 & s25_2;
process (clock_c) begin
  if rising_edge(clock_c) then
    if i5 = "1" then
      n3 <= "0";
    elsif i4 = "1" then
      n3 <= s29_2;
    end if;
  end if;
end process;
process (clock_c) begin
  if rising_edge(clock_c) then
    if i5 = "1" then
      n4 <= "0";
    elsif i4 = "1" then
      n4 <= n3;
    end if;
  end if;
end process;
process (clock_c) begin
  if rising_edge(clock_c) then
    if i5 = "1" then
      n5 <= "0";
    elsif i4 = "1" then
      n5 <= n4;
    end if;
  end if;
end process;
process (clock_c) begin
  if rising_edge(clock_c) then
    if i5 = "1" then
      n6 <= "0";
    elsif i4 = "1" then
      n6 <= n5;
    end if;
  end if;
end process;
n7 <= s29_1(10 downto 10) &
  s29_1(9 downto 9) &
  s29_1(8 downto 8) &
  s29_1(7 downto 7) &
  s29_1(6 downto 6) &
  s29_1(5 downto 5) &
  s29_1(4 downto 4) &
  s29_1(3 downto 3) &
  s29_1(2 downto 2) &
  s29_1(1 downto 1);
process (clock_c) begin
  if rising_edge(clock_c) then
    if i5 = "1" then
      n8 <= "0000000000";
    elsif i4 = "1" then
      n8 <= n7;
    end if;
  end if;
end process;
process (clock_c) begin
  if rising_edge(clock_c) then
    if i5 = "1" then
      n9 <= "0000000000";
    elsif i4 = "1" then
      n9 <= n8;
    end if;
  end if;
end process;
process (clock_c) begin
  if rising_edge(clock_c) then
    if i5 = "1" then
      n10 <= "0000000000";
    elsif i4 = "1" then
      n10 <= n9;
    end if;
  end if;
end process;
process (clock_c) begin
  if rising_edge(clock_c) then
    if i5 = "1" then
      n11 <= "0000000000";
    elsif i4 = "1" then
      n11 <= n10;
    end if;
  end if;
end process;
n12 <= s29_1(0 downto 0);
process (clock_c) begin
  if rising_edge(clock_c) then
    if i5 = "1" then
      n13 <= "0";
    elsif i4 = "1" then
      n13 <= n12;
    end if;
  end if;
end process;
process (clock_c) begin
  if rising_edge(clock_c) then
    if i5 = "1" then
      n14 <= "0";
    elsif i4 = "1" then
      n14 <= n13;
    end if;
  end if;
end process;
process (clock_c) begin
  if rising_edge(clock_c) then
    if i5 = "1" then
      n15 <= "0";
    elsif i4 = "1" then
      n15 <= n14;
    end if;
  end if;
end process;
process (clock_c) begin
  if rising_edge(clock_c) then
    if i5 = "1" then
      n16 <= "0";
    elsif i4 = "1" then
      n16 <= n15;
    end if;
  end if;
end process;
n17 <= not n16;
n18 <= s28_2 & s28_1;
n19 <= s28_3(71 downto 71) &
  s28_3(70 downto 70) &
  s28_3(69 downto 69) &
  s28_3(68 downto 68) &
  s28_3(67 downto 67) &
  s28_3(66 downto 66) &
  s28_3(65 downto 65) &
  s28_3(64 downto 64) &
  s28_3(63 downto 63) &
  s28_3(62 downto 62) &
  s28_3(61 downto 61) &
  s28_3(60 downto 60) &
  s28_3(59 downto 59) &
  s28_3(58 downto 58) &
  s28_3(57 downto 57) &
  s28_3(56 downto 56) &
  s28_3(55 downto 55) &
  s28_3(54 downto 54) &
  s28_3(53 downto 53) &
  s28_3(52 downto 52) &
  s28_3(51 downto 51) &
  s28_3(50 downto 50) &
  s28_3(49 downto 49) &
  s28_3(48 downto 48) &
  s28_3(47 downto 47) &
  s28_3(46 downto 46) &
  s28_3(45 downto 45) &
  s28_3(44 downto 44) &
  s28_3(43 downto 43) &
  s28_3(42 downto 42) &
  s28_3(41 downto 41) &
  s28_3(40 downto 40) &
  s28_3(39 downto 39) &
  s28_3(38 downto 38) &
  s28_3(37 downto 37) &
  s28_3(36 downto 36);
n20 <= s28_3(35 downto 35) &
  s28_3(34 downto 34) &
  s28_3(33 downto 33) &
  s28_3(32 downto 32) &
  s28_3(31 downto 31) &
  s28_3(30 downto 30) &
  s28_3(29 downto 29) &
  s28_3(28 downto 28) &
  s28_3(27 downto 27) &
  s28_3(26 downto 26) &
  s28_3(25 downto 25) &
  s28_3(24 downto 24) &
  s28_3(23 downto 23) &
  s28_3(22 downto 22) &
  s28_3(21 downto 21) &
  s28_3(20 downto 20) &
  s28_3(19 downto 19) &
  s28_3(18 downto 18) &
  s28_3(17 downto 17) &
  s28_3(16 downto 16) &
  s28_3(15 downto 15) &
  s28_3(14 downto 14) &
  s28_3(13 downto 13) &
  s28_3(12 downto 12) &
  s28_3(11 downto 11) &
  s28_3(10 downto 10) &
  s28_3(9 downto 9) &
  s28_3(8 downto 8) &
  s28_3(7 downto 7) &
  s28_3(6 downto 6) &
  s28_3(5 downto 5) &
  s28_3(4 downto 4) &
  s28_3(3 downto 3) &
  s28_3(2 downto 2) &
  s28_3(1 downto 1) &
  s28_3(0 downto 0);
n21 <= s27_1(71 downto 71) &
  s27_1(70 downto 70) &
  s27_1(69 downto 69) &
  s27_1(68 downto 68) &
  s27_1(67 downto 67) &
  s27_1(66 downto 66) &
  s27_1(65 downto 65) &
  s27_1(64 downto 64) &
  s27_1(63 downto 63) &
  s27_1(62 downto 62) &
  s27_1(61 downto 61) &
  s27_1(60 downto 60) &
  s27_1(59 downto 59) &
  s27_1(58 downto 58) &
  s27_1(57 downto 57) &
  s27_1(56 downto 56) &
  s27_1(55 downto 55) &
  s27_1(54 downto 54) &
  s27_1(53 downto 53) &
  s27_1(52 downto 52) &
  s27_1(51 downto 51) &
  s27_1(50 downto 50) &
  s27_1(49 downto 49) &
  s27_1(48 downto 48) &
  s27_1(47 downto 47) &
  s27_1(46 downto 46) &
  s27_1(45 downto 45) &
  s27_1(44 downto 44) &
  s27_1(43 downto 43) &
  s27_1(42 downto 42) &
  s27_1(41 downto 41) &
  s27_1(40 downto 40) &
  s27_1(39 downto 39) &
  s27_1(38 downto 38) &
  s27_1(37 downto 37) &
  s27_1(36 downto 36);
n22 <= s27_1(35 downto 35) &
  s27_1(34 downto 34) &
  s27_1(33 downto 33) &
  s27_1(32 downto 32) &
  s27_1(31 downto 31) &
  s27_1(30 downto 30) &
  s27_1(29 downto 29) &
  s27_1(28 downto 28) &
  s27_1(27 downto 27) &
  s27_1(26 downto 26) &
  s27_1(25 downto 25) &
  s27_1(24 downto 24) &
  s27_1(23 downto 23) &
  s27_1(22 downto 22) &
  s27_1(21 downto 21) &
  s27_1(20 downto 20) &
  s27_1(19 downto 19) &
  s27_1(18 downto 18) &
  s27_1(17 downto 17) &
  s27_1(16 downto 16) &
  s27_1(15 downto 15) &
  s27_1(14 downto 14) &
  s27_1(13 downto 13) &
  s27_1(12 downto 12) &
  s27_1(11 downto 11) &
  s27_1(10 downto 10) &
  s27_1(9 downto 9) &
  s27_1(8 downto 8) &
  s27_1(7 downto 7) &
  s27_1(6 downto 6) &
  s27_1(5 downto 5) &
  s27_1(4 downto 4) &
  s27_1(3 downto 3) &
  s27_1(2 downto 2) &
  s27_1(1 downto 1) &
  s27_1(0 downto 0);
n23 <= n20 when s26_1 = "1" else n19;
n24 <= n22 when s26_1 = "1" else n21;
s25 : cf_fft_4096_18_9 port map (clock_c, i2, i3, n1, i4, i5, s25_1, s25_2);
s26 : cf_fft_4096_18_37 port map (clock_c, n18, i4, i5, s26_1);
s27 : cf_fft_4096_18_33 port map (clock_c, n2, n6, n11, n16, i4, i5, s27_1);
s28 : cf_fft_4096_18_32 port map (clock_c, n2, n6, n11, n17, i4, i5, s28_1, s28_2, s28_3);
s29 : cf_fft_4096_18_28 port map (clock_c, i1, i4, i5, s29_1, s29_2);
o3 <= n24;
o2 <= n23;
o1 <= s28_1;
end architecture rtl;

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
entity cf_fft_4096_18_7 is
port (
clock_c : in std_logic;
i1 : in  unsigned(35 downto 0);
i2 : in  unsigned(35 downto 0);
i3 : in  unsigned(0 downto 0);
i4 : in  unsigned(0 downto 0);
i5 : in  unsigned(0 downto 0);
o1 : out unsigned(35 downto 0);
o2 : out unsigned(35 downto 0));
end entity cf_fft_4096_18_7;
architecture rtl of cf_fft_4096_18_7 is
signal n1 : unsigned(35 downto 0) := "000000000000000000000000000000000000";
signal n2 : unsigned(17 downto 0);
signal n3 : unsigned(17 downto 0);
signal n4 : unsigned(35 downto 0) := "000000000000000000000000000000000000";
signal n5 : unsigned(17 downto 0);
signal n6 : unsigned(17 downto 0);
signal n7 : unsigned(17 downto 0) := "000000000000000000";
signal n8 : unsigned(17 downto 0) := "000000000000000000";
signal n9 : unsigned(17 downto 0) := "000000000000000000";
signal n10 : unsigned(17 downto 0) := "000000000000000000";
signal n11 : unsigned(35 downto 0) := "000000000000000000000000000000000000";
signal n12 : unsigned(17 downto 0);
signal n13 : unsigned(17 downto 0);
signal n14 : unsigned(35 downto 0);
signal n15 : unsigned(17 downto 0);
signal n16 : unsigned(17 downto 0) := "000000000000000000";
signal n17 : unsigned(35 downto 0);
signal n18 : unsigned(17 downto 0);
signal n19 : unsigned(17 downto 0) := "000000000000000000";
signal n20 : unsigned(17 downto 0);
signal n21 : unsigned(17 downto 0) := "000000000000000000";
signal n22 : unsigned(35 downto 0);
signal n23 : unsigned(17 downto 0);
signal n24 : unsigned(17 downto 0) := "000000000000000000";
signal n25 : unsigned(35 downto 0);
signal n26 : unsigned(17 downto 0);
signal n27 : unsigned(17 downto 0) := "000000000000000000";
signal n28 : unsigned(17 downto 0);
signal n29 : unsigned(17 downto 0) := "000000000000000000";
signal n30 : unsigned(17 downto 0);
signal n31 : unsigned(17 downto 0);
signal n32 : unsigned(35 downto 0);
signal n33 : unsigned(35 downto 0) := "000000000000000000000000000000000000";
signal n34 : unsigned(17 downto 0);
signal n35 : unsigned(17 downto 0);
signal n36 : unsigned(35 downto 0);
signal n37 : unsigned(35 downto 0) := "000000000000000000000000000000000000";
begin
process (clock_c) begin
  if rising_edge(clock_c) then
    if i5 = "1" then
      n1 <= "000000000000000000000000000000000000";
    elsif i4 = "1" then
      n1 <= i1;
    end if;
  end if;
end process;
n2 <= n1(35 downto 35) &
  n1(34 downto 34) &
  n1(33 downto 33) &
  n1(32 downto 32) &
  n1(31 downto 31) &
  n1(30 downto 30) &
  n1(29 downto 29) &
  n1(28 downto 28) &
  n1(27 downto 27) &
  n1(26 downto 26) &
  n1(25 downto 25) &
  n1(24 downto 24) &
  n1(23 downto 23) &
  n1(22 downto 22) &
  n1(21 downto 21) &
  n1(20 downto 20) &
  n1(19 downto 19) &
  n1(18 downto 18);
n3 <= n1(17 downto 17) &
  n1(16 downto 16) &
  n1(15 downto 15) &
  n1(14 downto 14) &
  n1(13 downto 13) &
  n1(12 downto 12) &
  n1(11 downto 11) &
  n1(10 downto 10) &
  n1(9 downto 9) &
  n1(8 downto 8) &
  n1(7 downto 7) &
  n1(6 downto 6) &
  n1(5 downto 5) &
  n1(4 downto 4) &
  n1(3 downto 3) &
  n1(2 downto 2) &
  n1(1 downto 1) &
  n1(0 downto 0);
process (clock_c) begin
  if rising_edge(clock_c) then
    if i5 = "1" then
      n4 <= "000000000000000000000000000000000000";
    elsif i4 = "1" then
      n4 <= i2;
    end if;
  end if;
end process;
n5 <= n4(35 downto 35) &
  n4(34 downto 34) &
  n4(33 downto 33) &
  n4(32 downto 32) &
  n4(31 downto 31) &
  n4(30 downto 30) &
  n4(29 downto 29) &
  n4(28 downto 28) &
  n4(27 downto 27) &
  n4(26 downto 26) &
  n4(25 downto 25) &
  n4(24 downto 24) &
  n4(23 downto 23) &
  n4(22 downto 22) &
  n4(21 downto 21) &
  n4(20 downto 20) &
  n4(19 downto 19) &
  n4(18 downto 18);
n6 <= n4(17 downto 17) &
  n4(16 downto 16) &
  n4(15 downto 15) &
  n4(14 downto 14) &
  n4(13 downto 13) &
  n4(12 downto 12) &
  n4(11 downto 11) &
  n4(10 downto 10) &
  n4(9 downto 9) &
  n4(8 downto 8) &
  n4(7 downto 7) &
  n4(6 downto 6) &
  n4(5 downto 5) &
  n4(4 downto 4) &
  n4(3 downto 3) &
  n4(2 downto 2) &
  n4(1 downto 1) &
  n4(0 downto 0);
process (clock_c) begin
  if rising_edge(clock_c) then
    if i5 = "1" then
      n7 <= "000000000000000000";
    elsif i4 = "1" then
      n7 <= n2;
    end if;
  end if;
end process;
process (clock_c) begin
  if rising_edge(clock_c) then
    if i5 = "1" then
      n8 <= "000000000000000000";
    elsif i4 = "1" then
      n8 <= n7;
    end if;
  end if;
end process;
process (clock_c) begin
  if rising_edge(clock_c) then
    if i5 = "1" then
      n9 <= "000000000000000000";
    elsif i4 = "1" then
      n9 <= n3;
    end if;
  end if;
end process;
process (clock_c) begin
  if rising_edge(clock_c) then
    if i5 = "1" then
      n10 <= "000000000000000000";
    elsif i4 = "1" then
      n10 <= n9;
    end if;
  end if;
end process;
process (clock_c) begin
  if rising_edge(clock_c) then 
    if i4 = "1" then
      case i3 is
        when "0" => n11 <= "011111111111111111000000000000000000";
        when "1" => n11 <= "000000000000000000100000000000000000";
        when others => n11 <= "XXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX";
      end case;
    end if;
  end if;
end process;
n12 <= n11(35 downto 35) &
  n11(34 downto 34) &
  n11(33 downto 33) &
  n11(32 downto 32) &
  n11(31 downto 31) &
  n11(30 downto 30) &
  n11(29 downto 29) &
  n11(28 downto 28) &
  n11(27 downto 27) &
  n11(26 downto 26) &
  n11(25 downto 25) &
  n11(24 downto 24) &
  n11(23 downto 23) &
  n11(22 downto 22) &
  n11(21 downto 21) &
  n11(20 downto 20) &
  n11(19 downto 19) &
  n11(18 downto 18);
n13 <= n11(17 downto 17) &
  n11(16 downto 16) &
  n11(15 downto 15) &
  n11(14 downto 14) &
  n11(13 downto 13) &
  n11(12 downto 12) &
  n11(11 downto 11) &
  n11(10 downto 10) &
  n11(9 downto 9) &
  n11(8 downto 8) &
  n11(7 downto 7) &
  n11(6 downto 6) &
  n11(5 downto 5) &
  n11(4 downto 4) &
  n11(3 downto 3) &
  n11(2 downto 2) &
  n11(1 downto 1) &
  n11(0 downto 0);
n14 <= unsigned(signed(n5) * signed(n12));
n15 <= n14(34 downto 34) &
  n14(33 downto 33) &
  n14(32 downto 32) &
  n14(31 downto 31) &
  n14(30 downto 30) &
  n14(29 downto 29) &
  n14(28 downto 28) &
  n14(27 downto 27) &
  n14(26 downto 26) &
  n14(25 downto 25) &
  n14(24 downto 24) &
  n14(23 downto 23) &
  n14(22 downto 22) &
  n14(21 downto 21) &
  n14(20 downto 20) &
  n14(19 downto 19) &
  n14(18 downto 18) &
  n14(17 downto 17);
process (clock_c) begin
  if rising_edge(clock_c) then
    if i5 = "1" then
      n16 <= "000000000000000000";
    elsif i4 = "1" then
      n16 <= n15;
    end if;
  end if;
end process;
n17 <= unsigned(signed(n6) * signed(n13));
n18 <= n17(34 downto 34) &
  n17(33 downto 33) &
  n17(32 downto 32) &
  n17(31 downto 31) &
  n17(30 downto 30) &
  n17(29 downto 29) &
  n17(28 downto 28) &
  n17(27 downto 27) &
  n17(26 downto 26) &
  n17(25 downto 25) &
  n17(24 downto 24) &
  n17(23 downto 23) &
  n17(22 downto 22) &
  n17(21 downto 21) &
  n17(20 downto 20) &
  n17(19 downto 19) &
  n17(18 downto 18) &
  n17(17 downto 17);
process (clock_c) begin
  if rising_edge(clock_c) then
    if i5 = "1" then
      n19 <= "000000000000000000";
    elsif i4 = "1" then
      n19 <= n18;
    end if;
  end if;
end process;
n20 <= n16 - n19;
process (clock_c) begin
  if rising_edge(clock_c) then
    if i5 = "1" then
      n21 <= "000000000000000000";
    elsif i4 = "1" then
      n21 <= n20;
    end if;
  end if;
end process;
n22 <= unsigned(signed(n5) * signed(n13));
n23 <= n22(34 downto 34) &
  n22(33 downto 33) &
  n22(32 downto 32) &
  n22(31 downto 31) &
  n22(30 downto 30) &
  n22(29 downto 29) &
  n22(28 downto 28) &
  n22(27 downto 27) &
  n22(26 downto 26) &
  n22(25 downto 25) &
  n22(24 downto 24) &
  n22(23 downto 23) &
  n22(22 downto 22) &
  n22(21 downto 21) &
  n22(20 downto 20) &
  n22(19 downto 19) &
  n22(18 downto 18) &
  n22(17 downto 17);
process (clock_c) begin
  if rising_edge(clock_c) then
    if i5 = "1" then
      n24 <= "000000000000000000";
    elsif i4 = "1" then
      n24 <= n23;
    end if;
  end if;
end process;
n25 <= unsigned(signed(n6) * signed(n12));
n26 <= n25(34 downto 34) &
  n25(33 downto 33) &
  n25(32 downto 32) &
  n25(31 downto 31) &
  n25(30 downto 30) &
  n25(29 downto 29) &
  n25(28 downto 28) &
  n25(27 downto 27) &
  n25(26 downto 26) &
  n25(25 downto 25) &
  n25(24 downto 24) &
  n25(23 downto 23) &
  n25(22 downto 22) &
  n25(21 downto 21) &
  n25(20 downto 20) &
  n25(19 downto 19) &
  n25(18 downto 18) &
  n25(17 downto 17);
process (clock_c) begin
  if rising_edge(clock_c) then
    if i5 = "1" then
      n27 <= "000000000000000000";
    elsif i4 = "1" then
      n27 <= n26;
    end if;
  end if;
end process;
n28 <= n24 + n27;
process (clock_c) begin
  if rising_edge(clock_c) then
    if i5 = "1" then
      n29 <= "000000000000000000";
    elsif i4 = "1" then
      n29 <= n28;
    end if;
  end if;
end process;
n30 <= n8 + n21;
n31 <= n10 + n29;
n32 <= n30 & n31;
process (clock_c) begin
  if rising_edge(clock_c) then
    if i5 = "1" then
      n33 <= "000000000000000000000000000000000000";
    elsif i4 = "1" then
      n33 <= n32;
    end if;
  end if;
end process;
n34 <= n8 - n21;
n35 <= n10 - n29;
n36 <= n34 & n35;
process (clock_c) begin
  if rising_edge(clock_c) then
    if i5 = "1" then
      n37 <= "000000000000000000000000000000000000";
    elsif i4 = "1" then
      n37 <= n36;
    end if;
  end if;
end process;
o2 <= n37;
o1 <= n33;
end architecture rtl;

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
entity cf_fft_4096_18_6 is
port (
clock_c : in std_logic;
i1 : in  unsigned(0 downto 0);
i2 : in  unsigned(35 downto 0);
i3 : in  unsigned(35 downto 0);
i4 : in  unsigned(0 downto 0);
i5 : in  unsigned(0 downto 0);
o1 : out unsigned(0 downto 0);
o2 : out unsigned(35 downto 0);
o3 : out unsigned(35 downto 0));
end entity cf_fft_4096_18_6;
architecture rtl of cf_fft_4096_18_6 is
signal n1 : unsigned(0 downto 0);
signal n2 : unsigned(71 downto 0);
signal n3 : unsigned(0 downto 0) := "0";
signal n4 : unsigned(0 downto 0) := "0";
signal n5 : unsigned(0 downto 0) := "0";
signal n6 : unsigned(0 downto 0) := "0";
signal n7 : unsigned(9 downto 0);
signal n8 : unsigned(9 downto 0) := "0000000000";
signal n9 : unsigned(9 downto 0) := "0000000000";
signal n10 : unsigned(9 downto 0) := "0000000000";
signal n11 : unsigned(9 downto 0) := "0000000000";
signal n12 : unsigned(0 downto 0);
signal n13 : unsigned(0 downto 0) := "0";
signal n14 : unsigned(0 downto 0) := "0";
signal n15 : unsigned(0 downto 0) := "0";
signal n16 : unsigned(0 downto 0) := "0";
signal n17 : unsigned(0 downto 0);
signal n18 : unsigned(1 downto 0);
signal n19 : unsigned(35 downto 0);
signal n20 : unsigned(35 downto 0);
signal n21 : unsigned(35 downto 0);
signal n22 : unsigned(35 downto 0);
signal n23 : unsigned(35 downto 0);
signal n24 : unsigned(35 downto 0);
signal s25_1 : unsigned(35 downto 0);
signal s25_2 : unsigned(35 downto 0);
signal s26_1 : unsigned(0 downto 0);
signal s27_1 : unsigned(71 downto 0);
signal s28_1 : unsigned(0 downto 0);
signal s28_2 : unsigned(0 downto 0);
signal s28_3 : unsigned(71 downto 0);
signal s29_1 : unsigned(10 downto 0);
signal s29_2 : unsigned(0 downto 0);
component cf_fft_4096_18_7 is
port (
clock_c : in std_logic;
i1 : in  unsigned(35 downto 0);
i2 : in  unsigned(35 downto 0);
i3 : in  unsigned(0 downto 0);
i4 : in  unsigned(0 downto 0);
i5 : in  unsigned(0 downto 0);
o1 : out unsigned(35 downto 0);
o2 : out unsigned(35 downto 0));
end component cf_fft_4096_18_7;
component cf_fft_4096_18_37 is
port (
clock_c : in std_logic;
i1 : in  unsigned(1 downto 0);
i2 : in  unsigned(0 downto 0);
i3 : in  unsigned(0 downto 0);
o1 : out unsigned(0 downto 0));
end component cf_fft_4096_18_37;
component cf_fft_4096_18_33 is
port (
clock_c : in std_logic;
i1 : in  unsigned(71 downto 0);
i2 : in  unsigned(0 downto 0);
i3 : in  unsigned(9 downto 0);
i4 : in  unsigned(0 downto 0);
i5 : in  unsigned(0 downto 0);
i6 : in  unsigned(0 downto 0);
o1 : out unsigned(71 downto 0));
end component cf_fft_4096_18_33;
component cf_fft_4096_18_32 is
port (
clock_c : in std_logic;
i1 : in  unsigned(71 downto 0);
i2 : in  unsigned(0 downto 0);
i3 : in  unsigned(9 downto 0);
i4 : in  unsigned(0 downto 0);
i5 : in  unsigned(0 downto 0);
i6 : in  unsigned(0 downto 0);
o1 : out unsigned(0 downto 0);
o2 : out unsigned(0 downto 0);
o3 : out unsigned(71 downto 0));
end component cf_fft_4096_18_32;
component cf_fft_4096_18_28 is
port (
clock_c : in std_logic;
i1 : in  unsigned(0 downto 0);
i2 : in  unsigned(0 downto 0);
i3 : in  unsigned(0 downto 0);
o1 : out unsigned(10 downto 0);
o2 : out unsigned(0 downto 0));
end component cf_fft_4096_18_28;
begin
n1 <= s29_1(10 downto 10);
n2 <= s25_1 & s25_2;
process (clock_c) begin
  if rising_edge(clock_c) then
    if i5 = "1" then
      n3 <= "0";
    elsif i4 = "1" then
      n3 <= s29_2;
    end if;
  end if;
end process;
process (clock_c) begin
  if rising_edge(clock_c) then
    if i5 = "1" then
      n4 <= "0";
    elsif i4 = "1" then
      n4 <= n3;
    end if;
  end if;
end process;
process (clock_c) begin
  if rising_edge(clock_c) then
    if i5 = "1" then
      n5 <= "0";
    elsif i4 = "1" then
      n5 <= n4;
    end if;
  end if;
end process;
process (clock_c) begin
  if rising_edge(clock_c) then
    if i5 = "1" then
      n6 <= "0";
    elsif i4 = "1" then
      n6 <= n5;
    end if;
  end if;
end process;
n7 <= s29_1(10 downto 10) &
  s29_1(9 downto 9) &
  s29_1(8 downto 8) &
  s29_1(7 downto 7) &
  s29_1(6 downto 6) &
  s29_1(5 downto 5) &
  s29_1(4 downto 4) &
  s29_1(3 downto 3) &
  s29_1(2 downto 2) &
  s29_1(1 downto 1);
process (clock_c) begin
  if rising_edge(clock_c) then
    if i5 = "1" then
      n8 <= "0000000000";
    elsif i4 = "1" then
      n8 <= n7;
    end if;
  end if;
end process;
process (clock_c) begin
  if rising_edge(clock_c) then
    if i5 = "1" then
      n9 <= "0000000000";
    elsif i4 = "1" then
      n9 <= n8;
    end if;
  end if;
end process;
process (clock_c) begin
  if rising_edge(clock_c) then
    if i5 = "1" then
      n10 <= "0000000000";
    elsif i4 = "1" then
      n10 <= n9;
    end if;
  end if;
end process;
process (clock_c) begin
  if rising_edge(clock_c) then
    if i5 = "1" then
      n11 <= "0000000000";
    elsif i4 = "1" then
      n11 <= n10;
    end if;
  end if;
end process;
n12 <= s29_1(0 downto 0);
process (clock_c) begin
  if rising_edge(clock_c) then
    if i5 = "1" then
      n13 <= "0";
    elsif i4 = "1" then
      n13 <= n12;
    end if;
  end if;
end process;
process (clock_c) begin
  if rising_edge(clock_c) then
    if i5 = "1" then
      n14 <= "0";
    elsif i4 = "1" then
      n14 <= n13;
    end if;
  end if;
end process;
process (clock_c) begin
  if rising_edge(clock_c) then
    if i5 = "1" then
      n15 <= "0";
    elsif i4 = "1" then
      n15 <= n14;
    end if;
  end if;
end process;
process (clock_c) begin
  if rising_edge(clock_c) then
    if i5 = "1" then
      n16 <= "0";
    elsif i4 = "1" then
      n16 <= n15;
    end if;
  end if;
end process;
n17 <= not n16;
n18 <= s28_2 & s28_1;
n19 <= s28_3(71 downto 71) &
  s28_3(70 downto 70) &
  s28_3(69 downto 69) &
  s28_3(68 downto 68) &
  s28_3(67 downto 67) &
  s28_3(66 downto 66) &
  s28_3(65 downto 65) &
  s28_3(64 downto 64) &
  s28_3(63 downto 63) &
  s28_3(62 downto 62) &
  s28_3(61 downto 61) &
  s28_3(60 downto 60) &
  s28_3(59 downto 59) &
  s28_3(58 downto 58) &
  s28_3(57 downto 57) &
  s28_3(56 downto 56) &
  s28_3(55 downto 55) &
  s28_3(54 downto 54) &
  s28_3(53 downto 53) &
  s28_3(52 downto 52) &
  s28_3(51 downto 51) &
  s28_3(50 downto 50) &
  s28_3(49 downto 49) &
  s28_3(48 downto 48) &
  s28_3(47 downto 47) &
  s28_3(46 downto 46) &
  s28_3(45 downto 45) &
  s28_3(44 downto 44) &
  s28_3(43 downto 43) &
  s28_3(42 downto 42) &
  s28_3(41 downto 41) &
  s28_3(40 downto 40) &
  s28_3(39 downto 39) &
  s28_3(38 downto 38) &
  s28_3(37 downto 37) &
  s28_3(36 downto 36);
n20 <= s28_3(35 downto 35) &
  s28_3(34 downto 34) &
  s28_3(33 downto 33) &
  s28_3(32 downto 32) &
  s28_3(31 downto 31) &
  s28_3(30 downto 30) &
  s28_3(29 downto 29) &
  s28_3(28 downto 28) &
  s28_3(27 downto 27) &
  s28_3(26 downto 26) &
  s28_3(25 downto 25) &
  s28_3(24 downto 24) &
  s28_3(23 downto 23) &
  s28_3(22 downto 22) &
  s28_3(21 downto 21) &
  s28_3(20 downto 20) &
  s28_3(19 downto 19) &
  s28_3(18 downto 18) &
  s28_3(17 downto 17) &
  s28_3(16 downto 16) &
  s28_3(15 downto 15) &
  s28_3(14 downto 14) &
  s28_3(13 downto 13) &
  s28_3(12 downto 12) &
  s28_3(11 downto 11) &
  s28_3(10 downto 10) &
  s28_3(9 downto 9) &
  s28_3(8 downto 8) &
  s28_3(7 downto 7) &
  s28_3(6 downto 6) &
  s28_3(5 downto 5) &
  s28_3(4 downto 4) &
  s28_3(3 downto 3) &
  s28_3(2 downto 2) &
  s28_3(1 downto 1) &
  s28_3(0 downto 0);
n21 <= s27_1(71 downto 71) &
  s27_1(70 downto 70) &
  s27_1(69 downto 69) &
  s27_1(68 downto 68) &
  s27_1(67 downto 67) &
  s27_1(66 downto 66) &
  s27_1(65 downto 65) &
  s27_1(64 downto 64) &
  s27_1(63 downto 63) &
  s27_1(62 downto 62) &
  s27_1(61 downto 61) &
  s27_1(60 downto 60) &
  s27_1(59 downto 59) &
  s27_1(58 downto 58) &
  s27_1(57 downto 57) &
  s27_1(56 downto 56) &
  s27_1(55 downto 55) &
  s27_1(54 downto 54) &
  s27_1(53 downto 53) &
  s27_1(52 downto 52) &
  s27_1(51 downto 51) &
  s27_1(50 downto 50) &
  s27_1(49 downto 49) &
  s27_1(48 downto 48) &
  s27_1(47 downto 47) &
  s27_1(46 downto 46) &
  s27_1(45 downto 45) &
  s27_1(44 downto 44) &
  s27_1(43 downto 43) &
  s27_1(42 downto 42) &
  s27_1(41 downto 41) &
  s27_1(40 downto 40) &
  s27_1(39 downto 39) &
  s27_1(38 downto 38) &
  s27_1(37 downto 37) &
  s27_1(36 downto 36);
n22 <= s27_1(35 downto 35) &
  s27_1(34 downto 34) &
  s27_1(33 downto 33) &
  s27_1(32 downto 32) &
  s27_1(31 downto 31) &
  s27_1(30 downto 30) &
  s27_1(29 downto 29) &
  s27_1(28 downto 28) &
  s27_1(27 downto 27) &
  s27_1(26 downto 26) &
  s27_1(25 downto 25) &
  s27_1(24 downto 24) &
  s27_1(23 downto 23) &
  s27_1(22 downto 22) &
  s27_1(21 downto 21) &
  s27_1(20 downto 20) &
  s27_1(19 downto 19) &
  s27_1(18 downto 18) &
  s27_1(17 downto 17) &
  s27_1(16 downto 16) &
  s27_1(15 downto 15) &
  s27_1(14 downto 14) &
  s27_1(13 downto 13) &
  s27_1(12 downto 12) &
  s27_1(11 downto 11) &
  s27_1(10 downto 10) &
  s27_1(9 downto 9) &
  s27_1(8 downto 8) &
  s27_1(7 downto 7) &
  s27_1(6 downto 6) &
  s27_1(5 downto 5) &
  s27_1(4 downto 4) &
  s27_1(3 downto 3) &
  s27_1(2 downto 2) &
  s27_1(1 downto 1) &
  s27_1(0 downto 0);
n23 <= n20 when s26_1 = "1" else n19;
n24 <= n22 when s26_1 = "1" else n21;
s25 : cf_fft_4096_18_7 port map (clock_c, i2, i3, n1, i4, i5, s25_1, s25_2);
s26 : cf_fft_4096_18_37 port map (clock_c, n18, i4, i5, s26_1);
s27 : cf_fft_4096_18_33 port map (clock_c, n2, n6, n11, n16, i4, i5, s27_1);
s28 : cf_fft_4096_18_32 port map (clock_c, n2, n6, n11, n17, i4, i5, s28_1, s28_2, s28_3);
s29 : cf_fft_4096_18_28 port map (clock_c, i1, i4, i5, s29_1, s29_2);
o3 <= n24;
o2 <= n23;
o1 <= s28_1;
end architecture rtl;

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
entity cf_fft_4096_18_5 is
port (
clock_c : in std_logic;
i1 : in  unsigned(0 downto 0);
i2 : in  unsigned(35 downto 0);
i3 : in  unsigned(35 downto 0);
i4 : in  unsigned(0 downto 0);
i5 : in  unsigned(0 downto 0);
o1 : out unsigned(0 downto 0);
o2 : out unsigned(35 downto 0);
o3 : out unsigned(35 downto 0));
end entity cf_fft_4096_18_5;
architecture rtl of cf_fft_4096_18_5 is
signal n1 : unsigned(0 downto 0);
signal n2 : unsigned(71 downto 0);
signal n3 : unsigned(0 downto 0) := "0";
signal n4 : unsigned(0 downto 0) := "0";
signal n5 : unsigned(0 downto 0) := "0";
signal n6 : unsigned(0 downto 0) := "0";
signal n7 : unsigned(9 downto 0);
signal n8 : unsigned(9 downto 0) := "0000000000";
signal n9 : unsigned(9 downto 0) := "0000000000";
signal n10 : unsigned(9 downto 0) := "0000000000";
signal n11 : unsigned(9 downto 0) := "0000000000";
signal n12 : unsigned(0 downto 0);
signal n13 : unsigned(0 downto 0) := "0";
signal n14 : unsigned(0 downto 0) := "0";
signal n15 : unsigned(0 downto 0) := "0";
signal n16 : unsigned(0 downto 0) := "0";
signal n17 : unsigned(0 downto 0);
signal n18 : unsigned(1 downto 0);
signal n19 : unsigned(35 downto 0);
signal n20 : unsigned(35 downto 0);
signal n21 : unsigned(35 downto 0);
signal n22 : unsigned(35 downto 0);
signal n23 : unsigned(35 downto 0);
signal n24 : unsigned(35 downto 0);
signal s25_1 : unsigned(35 downto 0);
signal s25_2 : unsigned(35 downto 0);
signal s26_1 : unsigned(0 downto 0);
signal s27_1 : unsigned(71 downto 0);
signal s28_1 : unsigned(0 downto 0);
signal s28_2 : unsigned(0 downto 0);
signal s28_3 : unsigned(71 downto 0);
signal s29_1 : unsigned(10 downto 0);
signal s29_2 : unsigned(0 downto 0);
component cf_fft_4096_18_7 is
port (
clock_c : in std_logic;
i1 : in  unsigned(35 downto 0);
i2 : in  unsigned(35 downto 0);
i3 : in  unsigned(0 downto 0);
i4 : in  unsigned(0 downto 0);
i5 : in  unsigned(0 downto 0);
o1 : out unsigned(35 downto 0);
o2 : out unsigned(35 downto 0));
end component cf_fft_4096_18_7;
component cf_fft_4096_18_37 is
port (
clock_c : in std_logic;
i1 : in  unsigned(1 downto 0);
i2 : in  unsigned(0 downto 0);
i3 : in  unsigned(0 downto 0);
o1 : out unsigned(0 downto 0));
end component cf_fft_4096_18_37;
component cf_fft_4096_18_33 is
port (
clock_c : in std_logic;
i1 : in  unsigned(71 downto 0);
i2 : in  unsigned(0 downto 0);
i3 : in  unsigned(9 downto 0);
i4 : in  unsigned(0 downto 0);
i5 : in  unsigned(0 downto 0);
i6 : in  unsigned(0 downto 0);
o1 : out unsigned(71 downto 0));
end component cf_fft_4096_18_33;
component cf_fft_4096_18_32 is
port (
clock_c : in std_logic;
i1 : in  unsigned(71 downto 0);
i2 : in  unsigned(0 downto 0);
i3 : in  unsigned(9 downto 0);
i4 : in  unsigned(0 downto 0);
i5 : in  unsigned(0 downto 0);
i6 : in  unsigned(0 downto 0);
o1 : out unsigned(0 downto 0);
o2 : out unsigned(0 downto 0);
o3 : out unsigned(71 downto 0));
end component cf_fft_4096_18_32;
component cf_fft_4096_18_28 is
port (
clock_c : in std_logic;
i1 : in  unsigned(0 downto 0);
i2 : in  unsigned(0 downto 0);
i3 : in  unsigned(0 downto 0);
o1 : out unsigned(10 downto 0);
o2 : out unsigned(0 downto 0));
end component cf_fft_4096_18_28;
begin
n1 <= "0";
n2 <= s25_1 & s25_2;
process (clock_c) begin
  if rising_edge(clock_c) then
    if i5 = "1" then
      n3 <= "0";
    elsif i4 = "1" then
      n3 <= s29_2;
    end if;
  end if;
end process;
process (clock_c) begin
  if rising_edge(clock_c) then
    if i5 = "1" then
      n4 <= "0";
    elsif i4 = "1" then
      n4 <= n3;
    end if;
  end if;
end process;
process (clock_c) begin
  if rising_edge(clock_c) then
    if i5 = "1" then
      n5 <= "0";
    elsif i4 = "1" then
      n5 <= n4;
    end if;
  end if;
end process;
process (clock_c) begin
  if rising_edge(clock_c) then
    if i5 = "1" then
      n6 <= "0";
    elsif i4 = "1" then
      n6 <= n5;
    end if;
  end if;
end process;
n7 <= s29_1(10 downto 10) &
  s29_1(9 downto 9) &
  s29_1(8 downto 8) &
  s29_1(7 downto 7) &
  s29_1(6 downto 6) &
  s29_1(5 downto 5) &
  s29_1(4 downto 4) &
  s29_1(3 downto 3) &
  s29_1(2 downto 2) &
  s29_1(1 downto 1);
process (clock_c) begin
  if rising_edge(clock_c) then
    if i5 = "1" then
      n8 <= "0000000000";
    elsif i4 = "1" then
      n8 <= n7;
    end if;
  end if;
end process;
process (clock_c) begin
  if rising_edge(clock_c) then
    if i5 = "1" then
      n9 <= "0000000000";
    elsif i4 = "1" then
      n9 <= n8;
    end if;
  end if;
end process;
process (clock_c) begin
  if rising_edge(clock_c) then
    if i5 = "1" then
      n10 <= "0000000000";
    elsif i4 = "1" then
      n10 <= n9;
    end if;
  end if;
end process;
process (clock_c) begin
  if rising_edge(clock_c) then
    if i5 = "1" then
      n11 <= "0000000000";
    elsif i4 = "1" then
      n11 <= n10;
    end if;
  end if;
end process;
n12 <= s29_1(0 downto 0);
process (clock_c) begin
  if rising_edge(clock_c) then
    if i5 = "1" then
      n13 <= "0";
    elsif i4 = "1" then
      n13 <= n12;
    end if;
  end if;
end process;
process (clock_c) begin
  if rising_edge(clock_c) then
    if i5 = "1" then
      n14 <= "0";
    elsif i4 = "1" then
      n14 <= n13;
    end if;
  end if;
end process;
process (clock_c) begin
  if rising_edge(clock_c) then
    if i5 = "1" then
      n15 <= "0";
    elsif i4 = "1" then
      n15 <= n14;
    end if;
  end if;
end process;
process (clock_c) begin
  if rising_edge(clock_c) then
    if i5 = "1" then
      n16 <= "0";
    elsif i4 = "1" then
      n16 <= n15;
    end if;
  end if;
end process;
n17 <= not n16;
n18 <= s28_2 & s28_1;
n19 <= s28_3(71 downto 71) &
  s28_3(70 downto 70) &
  s28_3(69 downto 69) &
  s28_3(68 downto 68) &
  s28_3(67 downto 67) &
  s28_3(66 downto 66) &
  s28_3(65 downto 65) &
  s28_3(64 downto 64) &
  s28_3(63 downto 63) &
  s28_3(62 downto 62) &
  s28_3(61 downto 61) &
  s28_3(60 downto 60) &
  s28_3(59 downto 59) &
  s28_3(58 downto 58) &
  s28_3(57 downto 57) &
  s28_3(56 downto 56) &
  s28_3(55 downto 55) &
  s28_3(54 downto 54) &
  s28_3(53 downto 53) &
  s28_3(52 downto 52) &
  s28_3(51 downto 51) &
  s28_3(50 downto 50) &
  s28_3(49 downto 49) &
  s28_3(48 downto 48) &
  s28_3(47 downto 47) &
  s28_3(46 downto 46) &
  s28_3(45 downto 45) &
  s28_3(44 downto 44) &
  s28_3(43 downto 43) &
  s28_3(42 downto 42) &
  s28_3(41 downto 41) &
  s28_3(40 downto 40) &
  s28_3(39 downto 39) &
  s28_3(38 downto 38) &
  s28_3(37 downto 37) &
  s28_3(36 downto 36);
n20 <= s28_3(35 downto 35) &
  s28_3(34 downto 34) &
  s28_3(33 downto 33) &
  s28_3(32 downto 32) &
  s28_3(31 downto 31) &
  s28_3(30 downto 30) &
  s28_3(29 downto 29) &
  s28_3(28 downto 28) &
  s28_3(27 downto 27) &
  s28_3(26 downto 26) &
  s28_3(25 downto 25) &
  s28_3(24 downto 24) &
  s28_3(23 downto 23) &
  s28_3(22 downto 22) &
  s28_3(21 downto 21) &
  s28_3(20 downto 20) &
  s28_3(19 downto 19) &
  s28_3(18 downto 18) &
  s28_3(17 downto 17) &
  s28_3(16 downto 16) &
  s28_3(15 downto 15) &
  s28_3(14 downto 14) &
  s28_3(13 downto 13) &
  s28_3(12 downto 12) &
  s28_3(11 downto 11) &
  s28_3(10 downto 10) &
  s28_3(9 downto 9) &
  s28_3(8 downto 8) &
  s28_3(7 downto 7) &
  s28_3(6 downto 6) &
  s28_3(5 downto 5) &
  s28_3(4 downto 4) &
  s28_3(3 downto 3) &
  s28_3(2 downto 2) &
  s28_3(1 downto 1) &
  s28_3(0 downto 0);
n21 <= s27_1(71 downto 71) &
  s27_1(70 downto 70) &
  s27_1(69 downto 69) &
  s27_1(68 downto 68) &
  s27_1(67 downto 67) &
  s27_1(66 downto 66) &
  s27_1(65 downto 65) &
  s27_1(64 downto 64) &
  s27_1(63 downto 63) &
  s27_1(62 downto 62) &
  s27_1(61 downto 61) &
  s27_1(60 downto 60) &
  s27_1(59 downto 59) &
  s27_1(58 downto 58) &
  s27_1(57 downto 57) &
  s27_1(56 downto 56) &
  s27_1(55 downto 55) &
  s27_1(54 downto 54) &
  s27_1(53 downto 53) &
  s27_1(52 downto 52) &
  s27_1(51 downto 51) &
  s27_1(50 downto 50) &
  s27_1(49 downto 49) &
  s27_1(48 downto 48) &
  s27_1(47 downto 47) &
  s27_1(46 downto 46) &
  s27_1(45 downto 45) &
  s27_1(44 downto 44) &
  s27_1(43 downto 43) &
  s27_1(42 downto 42) &
  s27_1(41 downto 41) &
  s27_1(40 downto 40) &
  s27_1(39 downto 39) &
  s27_1(38 downto 38) &
  s27_1(37 downto 37) &
  s27_1(36 downto 36);
n22 <= s27_1(35 downto 35) &
  s27_1(34 downto 34) &
  s27_1(33 downto 33) &
  s27_1(32 downto 32) &
  s27_1(31 downto 31) &
  s27_1(30 downto 30) &
  s27_1(29 downto 29) &
  s27_1(28 downto 28) &
  s27_1(27 downto 27) &
  s27_1(26 downto 26) &
  s27_1(25 downto 25) &
  s27_1(24 downto 24) &
  s27_1(23 downto 23) &
  s27_1(22 downto 22) &
  s27_1(21 downto 21) &
  s27_1(20 downto 20) &
  s27_1(19 downto 19) &
  s27_1(18 downto 18) &
  s27_1(17 downto 17) &
  s27_1(16 downto 16) &
  s27_1(15 downto 15) &
  s27_1(14 downto 14) &
  s27_1(13 downto 13) &
  s27_1(12 downto 12) &
  s27_1(11 downto 11) &
  s27_1(10 downto 10) &
  s27_1(9 downto 9) &
  s27_1(8 downto 8) &
  s27_1(7 downto 7) &
  s27_1(6 downto 6) &
  s27_1(5 downto 5) &
  s27_1(4 downto 4) &
  s27_1(3 downto 3) &
  s27_1(2 downto 2) &
  s27_1(1 downto 1) &
  s27_1(0 downto 0);
n23 <= n20 when s26_1 = "1" else n19;
n24 <= n22 when s26_1 = "1" else n21;
s25 : cf_fft_4096_18_7 port map (clock_c, i2, i3, n1, i4, i5, s25_1, s25_2);
s26 : cf_fft_4096_18_37 port map (clock_c, n18, i4, i5, s26_1);
s27 : cf_fft_4096_18_33 port map (clock_c, n2, n6, n11, n16, i4, i5, s27_1);
s28 : cf_fft_4096_18_32 port map (clock_c, n2, n6, n11, n17, i4, i5, s28_1, s28_2, s28_3);
s29 : cf_fft_4096_18_28 port map (clock_c, i1, i4, i5, s29_1, s29_2);
o3 <= n24;
o2 <= n23;
o1 <= s28_1;
end architecture rtl;

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
entity cf_fft_4096_18_4 is
port (
clock_c : in std_logic;
i1 : in  unsigned(0 downto 0);
i2 : in  unsigned(71 downto 0);
i3 : in  unsigned(0 downto 0);
i4 : in  unsigned(9 downto 0);
i5 : in  unsigned(0 downto 0);
i6 : in  unsigned(0 downto 0);
o1 : out unsigned(71 downto 0));
end entity cf_fft_4096_18_4;
architecture rtl of cf_fft_4096_18_4 is
signal n1 : unsigned(9 downto 0);
signal n2 : unsigned(9 downto 0);
signal n3 : unsigned(9 downto 0) := "0000000000";
signal n4 : unsigned(0 downto 0);
signal n5 : unsigned(0 downto 0);
signal n6 : unsigned(71 downto 0);
signal n6a : unsigned(9 downto 0) := "0000000000";
type   n6mt is array (1023 downto 0) of unsigned(71 downto 0);
signal n6m : n6mt;
signal n7 : unsigned(0 downto 0);
signal n8 : unsigned(71 downto 0);
signal n8a : unsigned(9 downto 0) := "0000000000";
type   n8mt is array (1023 downto 0) of unsigned(71 downto 0);
signal n8m : n8mt;
signal n9 : unsigned(0 downto 0) := "0";
signal n10 : unsigned(71 downto 0);
signal n11 : unsigned(0 downto 0);
signal s12_1 : unsigned(0 downto 0);
component cf_fft_4096_18_34 is
port (
clock_c : in std_logic;
i1 : in  unsigned(0 downto 0);
i2 : in  unsigned(0 downto 0);
i3 : in  unsigned(0 downto 0);
o1 : out unsigned(0 downto 0));
end component cf_fft_4096_18_34;
begin
n1 <= "0000000001";
n2 <= n3 + n1;
process (clock_c) begin
  if rising_edge(clock_c) then
    if n11 = "1" then
      n3 <= "0000000000";
    elsif i5 = "1" then
      n3 <= n2;
    end if;
  end if;
end process;
n4 <= not s12_1;
n5 <= i3 and n4;
process (clock_c) begin
  if rising_edge(clock_c) then
    if i5 = "1" then
      if n5 = "1" then
        n6m(to_integer(i4)) <= i2;
      end if;
      n6a <= n3;
    end if;
  end if;
end process;
n6 <= n6m(to_integer(n6a));
n7 <= i3 and s12_1;
process (clock_c) begin
  if rising_edge(clock_c) then
    if i5 = "1" then
      if n7 = "1" then
        n8m(to_integer(i4)) <= i2;
      end if;
      n8a <= n3;
    end if;
  end if;
end process;
n8 <= n8m(to_integer(n8a));
process (clock_c) begin
  if rising_edge(clock_c) then
    if i6 = "1" then
      n9 <= "0";
    elsif i5 = "1" then
      n9 <= n4;
    end if;
  end if;
end process;
n10 <= n8 when n9 = "1" else n6;
n11 <= i1 or i6;
s12 : cf_fft_4096_18_34 port map (clock_c, i1, i5, i6, s12_1);
o1 <= n10;
end architecture rtl;

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
entity cf_fft_4096_18_3 is
port (
clock_c : in std_logic;
i1 : in  unsigned(0 downto 0);
i2 : in  unsigned(71 downto 0);
i3 : in  unsigned(0 downto 0);
i4 : in  unsigned(9 downto 0);
i5 : in  unsigned(0 downto 0);
i6 : in  unsigned(0 downto 0);
o1 : out unsigned(0 downto 0);
o2 : out unsigned(0 downto 0);
o3 : out unsigned(71 downto 0));
end entity cf_fft_4096_18_3;
architecture rtl of cf_fft_4096_18_3 is
signal n1 : unsigned(9 downto 0);
signal n2 : unsigned(9 downto 0);
signal n3 : unsigned(9 downto 0) := "0000000000";
signal n4 : unsigned(0 downto 0);
signal n5 : unsigned(0 downto 0) := "0";
signal n6 : unsigned(9 downto 0);
signal n7 : unsigned(0 downto 0);
signal n8 : unsigned(0 downto 0);
signal n9 : unsigned(71 downto 0);
signal n9a : unsigned(9 downto 0) := "0000000000";
type   n9mt is array (1023 downto 0) of unsigned(71 downto 0);
signal n9m : n9mt;
signal n10 : unsigned(0 downto 0);
signal n11 : unsigned(71 downto 0);
signal n11a : unsigned(9 downto 0) := "0000000000";
type   n11mt is array (1023 downto 0) of unsigned(71 downto 0);
signal n11m : n11mt;
signal n12 : unsigned(0 downto 0) := "0";
signal n13 : unsigned(71 downto 0);
signal n14 : unsigned(0 downto 0);
signal s15_1 : unsigned(0 downto 0);
component cf_fft_4096_18_34 is
port (
clock_c : in std_logic;
i1 : in  unsigned(0 downto 0);
i2 : in  unsigned(0 downto 0);
i3 : in  unsigned(0 downto 0);
o1 : out unsigned(0 downto 0));
end component cf_fft_4096_18_34;
begin
n1 <= "0000000001";
n2 <= n3 + n1;
process (clock_c) begin
  if rising_edge(clock_c) then
    if n14 = "1" then
      n3 <= "0000000000";
    elsif i5 = "1" then
      n3 <= n2;
    end if;
  end if;
end process;
n4 <= not s15_1;
process (clock_c) begin
  if rising_edge(clock_c) then
    if i6 = "1" then
      n5 <= "0";
    elsif i5 = "1" then
      n5 <= i1;
    end if;
  end if;
end process;
n6 <= "0000000000";
n7 <= "1" when n3 = n6 else "0";
n8 <= i3 and n4;
process (clock_c) begin
  if rising_edge(clock_c) then
    if i5 = "1" then
      if n8 = "1" then
        n9m(to_integer(i4)) <= i2;
      end if;
      n9a <= n3;
    end if;
  end if;
end process;
n9 <= n9m(to_integer(n9a));
n10 <= i3 and s15_1;
process (clock_c) begin
  if rising_edge(clock_c) then
    if i5 = "1" then
      if n10 = "1" then
        n11m(to_integer(i4)) <= i2;
      end if;
      n11a <= n3;
    end if;
  end if;
end process;
n11 <= n11m(to_integer(n11a));
process (clock_c) begin
  if rising_edge(clock_c) then
    if i6 = "1" then
      n12 <= "0";
    elsif i5 = "1" then
      n12 <= n4;
    end if;
  end if;
end process;
n13 <= n11 when n12 = "1" else n9;
n14 <= i1 or i6;
s15 : cf_fft_4096_18_34 port map (clock_c, i1, i5, i6, s15_1);
o3 <= n13;
o2 <= n7;
o1 <= n5;
end architecture rtl;

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
entity cf_fft_4096_18_2 is
port (
clock_c : in std_logic;
i1 : in  unsigned(0 downto 0);
i2 : in  unsigned(35 downto 0);
i3 : in  unsigned(35 downto 0);
i4 : in  unsigned(0 downto 0);
i5 : in  unsigned(0 downto 0);
o1 : out unsigned(0 downto 0);
o2 : out unsigned(35 downto 0);
o3 : out unsigned(35 downto 0));
end entity cf_fft_4096_18_2;
architecture rtl of cf_fft_4096_18_2 is
signal n1 : unsigned(71 downto 0);
signal n2 : unsigned(0 downto 0);
signal n3 : unsigned(0 downto 0);
signal n4 : unsigned(9 downto 0);
signal n5 : unsigned(9 downto 0);
signal n6 : unsigned(1 downto 0);
signal n7 : unsigned(35 downto 0);
signal n8 : unsigned(35 downto 0);
signal n9 : unsigned(35 downto 0);
signal n10 : unsigned(35 downto 0);
signal n11 : unsigned(35 downto 0);
signal n12 : unsigned(35 downto 0);
signal s13_1 : unsigned(0 downto 0);
signal s14_1 : unsigned(71 downto 0);
signal s15_1 : unsigned(0 downto 0);
signal s15_2 : unsigned(0 downto 0);
signal s15_3 : unsigned(71 downto 0);
signal s16_1 : unsigned(10 downto 0);
signal s16_2 : unsigned(0 downto 0);
component cf_fft_4096_18_37 is
port (
clock_c : in std_logic;
i1 : in  unsigned(1 downto 0);
i2 : in  unsigned(0 downto 0);
i3 : in  unsigned(0 downto 0);
o1 : out unsigned(0 downto 0));
end component cf_fft_4096_18_37;
component cf_fft_4096_18_4 is
port (
clock_c : in std_logic;
i1 : in  unsigned(0 downto 0);
i2 : in  unsigned(71 downto 0);
i3 : in  unsigned(0 downto 0);
i4 : in  unsigned(9 downto 0);
i5 : in  unsigned(0 downto 0);
i6 : in  unsigned(0 downto 0);
o1 : out unsigned(71 downto 0));
end component cf_fft_4096_18_4;
component cf_fft_4096_18_3 is
port (
clock_c : in std_logic;
i1 : in  unsigned(0 downto 0);
i2 : in  unsigned(71 downto 0);
i3 : in  unsigned(0 downto 0);
i4 : in  unsigned(9 downto 0);
i5 : in  unsigned(0 downto 0);
i6 : in  unsigned(0 downto 0);
o1 : out unsigned(0 downto 0);
o2 : out unsigned(0 downto 0);
o3 : out unsigned(71 downto 0));
end component cf_fft_4096_18_3;
component cf_fft_4096_18_28 is
port (
clock_c : in std_logic;
i1 : in  unsigned(0 downto 0);
i2 : in  unsigned(0 downto 0);
i3 : in  unsigned(0 downto 0);
o1 : out unsigned(10 downto 0);
o2 : out unsigned(0 downto 0));
end component cf_fft_4096_18_28;
begin
n1 <= i2 & i3;
n2 <= s16_1(10 downto 10);
n3 <= not n2;
n4 <= s16_1(9 downto 9) &
  s16_1(8 downto 8) &
  s16_1(7 downto 7) &
  s16_1(6 downto 6) &
  s16_1(5 downto 5) &
  s16_1(4 downto 4) &
  s16_1(3 downto 3) &
  s16_1(2 downto 2) &
  s16_1(1 downto 1) &
  s16_1(0 downto 0);
n5 <= n4(0 downto 0) &
  n4(1 downto 1) &
  n4(2 downto 2) &
  n4(3 downto 3) &
  n4(4 downto 4) &
  n4(5 downto 5) &
  n4(6 downto 6) &
  n4(7 downto 7) &
  n4(8 downto 8) &
  n4(9 downto 9);
n6 <= s15_2 & s15_1;
n7 <= s15_3(71 downto 71) &
  s15_3(70 downto 70) &
  s15_3(69 downto 69) &
  s15_3(68 downto 68) &
  s15_3(67 downto 67) &
  s15_3(66 downto 66) &
  s15_3(65 downto 65) &
  s15_3(64 downto 64) &
  s15_3(63 downto 63) &
  s15_3(62 downto 62) &
  s15_3(61 downto 61) &
  s15_3(60 downto 60) &
  s15_3(59 downto 59) &
  s15_3(58 downto 58) &
  s15_3(57 downto 57) &
  s15_3(56 downto 56) &
  s15_3(55 downto 55) &
  s15_3(54 downto 54) &
  s15_3(53 downto 53) &
  s15_3(52 downto 52) &
  s15_3(51 downto 51) &
  s15_3(50 downto 50) &
  s15_3(49 downto 49) &
  s15_3(48 downto 48) &
  s15_3(47 downto 47) &
  s15_3(46 downto 46) &
  s15_3(45 downto 45) &
  s15_3(44 downto 44) &
  s15_3(43 downto 43) &
  s15_3(42 downto 42) &
  s15_3(41 downto 41) &
  s15_3(40 downto 40) &
  s15_3(39 downto 39) &
  s15_3(38 downto 38) &
  s15_3(37 downto 37) &
  s15_3(36 downto 36);
n8 <= s15_3(35 downto 35) &
  s15_3(34 downto 34) &
  s15_3(33 downto 33) &
  s15_3(32 downto 32) &
  s15_3(31 downto 31) &
  s15_3(30 downto 30) &
  s15_3(29 downto 29) &
  s15_3(28 downto 28) &
  s15_3(27 downto 27) &
  s15_3(26 downto 26) &
  s15_3(25 downto 25) &
  s15_3(24 downto 24) &
  s15_3(23 downto 23) &
  s15_3(22 downto 22) &
  s15_3(21 downto 21) &
  s15_3(20 downto 20) &
  s15_3(19 downto 19) &
  s15_3(18 downto 18) &
  s15_3(17 downto 17) &
  s15_3(16 downto 16) &
  s15_3(15 downto 15) &
  s15_3(14 downto 14) &
  s15_3(13 downto 13) &
  s15_3(12 downto 12) &
  s15_3(11 downto 11) &
  s15_3(10 downto 10) &
  s15_3(9 downto 9) &
  s15_3(8 downto 8) &
  s15_3(7 downto 7) &
  s15_3(6 downto 6) &
  s15_3(5 downto 5) &
  s15_3(4 downto 4) &
  s15_3(3 downto 3) &
  s15_3(2 downto 2) &
  s15_3(1 downto 1) &
  s15_3(0 downto 0);
n9 <= s14_1(71 downto 71) &
  s14_1(70 downto 70) &
  s14_1(69 downto 69) &
  s14_1(68 downto 68) &
  s14_1(67 downto 67) &
  s14_1(66 downto 66) &
  s14_1(65 downto 65) &
  s14_1(64 downto 64) &
  s14_1(63 downto 63) &
  s14_1(62 downto 62) &
  s14_1(61 downto 61) &
  s14_1(60 downto 60) &
  s14_1(59 downto 59) &
  s14_1(58 downto 58) &
  s14_1(57 downto 57) &
  s14_1(56 downto 56) &
  s14_1(55 downto 55) &
  s14_1(54 downto 54) &
  s14_1(53 downto 53) &
  s14_1(52 downto 52) &
  s14_1(51 downto 51) &
  s14_1(50 downto 50) &
  s14_1(49 downto 49) &
  s14_1(48 downto 48) &
  s14_1(47 downto 47) &
  s14_1(46 downto 46) &
  s14_1(45 downto 45) &
  s14_1(44 downto 44) &
  s14_1(43 downto 43) &
  s14_1(42 downto 42) &
  s14_1(41 downto 41) &
  s14_1(40 downto 40) &
  s14_1(39 downto 39) &
  s14_1(38 downto 38) &
  s14_1(37 downto 37) &
  s14_1(36 downto 36);
n10 <= s14_1(35 downto 35) &
  s14_1(34 downto 34) &
  s14_1(33 downto 33) &
  s14_1(32 downto 32) &
  s14_1(31 downto 31) &
  s14_1(30 downto 30) &
  s14_1(29 downto 29) &
  s14_1(28 downto 28) &
  s14_1(27 downto 27) &
  s14_1(26 downto 26) &
  s14_1(25 downto 25) &
  s14_1(24 downto 24) &
  s14_1(23 downto 23) &
  s14_1(22 downto 22) &
  s14_1(21 downto 21) &
  s14_1(20 downto 20) &
  s14_1(19 downto 19) &
  s14_1(18 downto 18) &
  s14_1(17 downto 17) &
  s14_1(16 downto 16) &
  s14_1(15 downto 15) &
  s14_1(14 downto 14) &
  s14_1(13 downto 13) &
  s14_1(12 downto 12) &
  s14_1(11 downto 11) &
  s14_1(10 downto 10) &
  s14_1(9 downto 9) &
  s14_1(8 downto 8) &
  s14_1(7 downto 7) &
  s14_1(6 downto 6) &
  s14_1(5 downto 5) &
  s14_1(4 downto 4) &
  s14_1(3 downto 3) &
  s14_1(2 downto 2) &
  s14_1(1 downto 1) &
  s14_1(0 downto 0);
n11 <= n8 when s13_1 = "1" else n7;
n12 <= n10 when s13_1 = "1" else n9;
s13 : cf_fft_4096_18_37 port map (clock_c, n6, i4, i5, s13_1);
s14 : cf_fft_4096_18_4 port map (clock_c, s16_2, n1, n2, n5, i4, i5, s14_1);
s15 : cf_fft_4096_18_3 port map (clock_c, s16_2, n1, n3, n5, i4, i5, s15_1, s15_2, s15_3);
s16 : cf_fft_4096_18_28 port map (clock_c, i1, i4, i5, s16_1, s16_2);
o3 <= n12;
o2 <= n11;
o1 <= s15_1;
end architecture rtl;

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
entity cf_fft_4096_18_1 is
port (
clock_c : in std_logic;
i1 : in  unsigned(0 downto 0);
i2 : in  unsigned(35 downto 0);
i3 : in  unsigned(35 downto 0);
i4 : in  unsigned(0 downto 0);
i5 : in  unsigned(0 downto 0);
o1 : out unsigned(0 downto 0);
o2 : out unsigned(35 downto 0);
o3 : out unsigned(35 downto 0));
end entity cf_fft_4096_18_1;
architecture rtl of cf_fft_4096_18_1 is
signal s1_1 : unsigned(0 downto 0);
signal s1_2 : unsigned(35 downto 0);
signal s1_3 : unsigned(35 downto 0);
signal s2_1 : unsigned(0 downto 0);
signal s2_2 : unsigned(35 downto 0);
signal s2_3 : unsigned(35 downto 0);
signal s3_1 : unsigned(0 downto 0);
signal s3_2 : unsigned(35 downto 0);
signal s3_3 : unsigned(35 downto 0);
signal s4_1 : unsigned(0 downto 0);
signal s4_2 : unsigned(35 downto 0);
signal s4_3 : unsigned(35 downto 0);
signal s5_1 : unsigned(0 downto 0);
signal s5_2 : unsigned(35 downto 0);
signal s5_3 : unsigned(35 downto 0);
signal s6_1 : unsigned(0 downto 0);
signal s6_2 : unsigned(35 downto 0);
signal s6_3 : unsigned(35 downto 0);
component cf_fft_4096_18_27 is
port (
clock_c : in std_logic;
i1 : in  unsigned(0 downto 0);
i2 : in  unsigned(35 downto 0);
i3 : in  unsigned(35 downto 0);
i4 : in  unsigned(0 downto 0);
i5 : in  unsigned(0 downto 0);
o1 : out unsigned(0 downto 0);
o2 : out unsigned(35 downto 0);
o3 : out unsigned(35 downto 0));
end component cf_fft_4096_18_27;
component cf_fft_4096_18_10 is
port (
clock_c : in std_logic;
i1 : in  unsigned(0 downto 0);
i2 : in  unsigned(35 downto 0);
i3 : in  unsigned(35 downto 0);
i4 : in  unsigned(0 downto 0);
i5 : in  unsigned(0 downto 0);
o1 : out unsigned(0 downto 0);
o2 : out unsigned(35 downto 0);
o3 : out unsigned(35 downto 0));
end component cf_fft_4096_18_10;
component cf_fft_4096_18_8 is
port (
clock_c : in std_logic;
i1 : in  unsigned(0 downto 0);
i2 : in  unsigned(35 downto 0);
i3 : in  unsigned(35 downto 0);
i4 : in  unsigned(0 downto 0);
i5 : in  unsigned(0 downto 0);
o1 : out unsigned(0 downto 0);
o2 : out unsigned(35 downto 0);
o3 : out unsigned(35 downto 0));
end component cf_fft_4096_18_8;
component cf_fft_4096_18_6 is
port (
clock_c : in std_logic;
i1 : in  unsigned(0 downto 0);
i2 : in  unsigned(35 downto 0);
i3 : in  unsigned(35 downto 0);
i4 : in  unsigned(0 downto 0);
i5 : in  unsigned(0 downto 0);
o1 : out unsigned(0 downto 0);
o2 : out unsigned(35 downto 0);
o3 : out unsigned(35 downto 0));
end component cf_fft_4096_18_6;
component cf_fft_4096_18_5 is
port (
clock_c : in std_logic;
i1 : in  unsigned(0 downto 0);
i2 : in  unsigned(35 downto 0);
i3 : in  unsigned(35 downto 0);
i4 : in  unsigned(0 downto 0);
i5 : in  unsigned(0 downto 0);
o1 : out unsigned(0 downto 0);
o2 : out unsigned(35 downto 0);
o3 : out unsigned(35 downto 0));
end component cf_fft_4096_18_5;
component cf_fft_4096_18_2 is
port (
clock_c : in std_logic;
i1 : in  unsigned(0 downto 0);
i2 : in  unsigned(35 downto 0);
i3 : in  unsigned(35 downto 0);
i4 : in  unsigned(0 downto 0);
i5 : in  unsigned(0 downto 0);
o1 : out unsigned(0 downto 0);
o2 : out unsigned(35 downto 0);
o3 : out unsigned(35 downto 0));
end component cf_fft_4096_18_2;
begin
s1 : cf_fft_4096_18_27 port map (clock_c, s3_1, s3_2, s3_3, i4, i5, s1_1, s1_2, s1_3);
s2 : cf_fft_4096_18_10 port map (clock_c, s1_1, s1_2, s1_3, i4, i5, s2_1, s2_2, s2_3);
s3 : cf_fft_4096_18_8 port map (clock_c, s4_1, s4_2, s4_3, i4, i5, s3_1, s3_2, s3_3);
s4 : cf_fft_4096_18_6 port map (clock_c, s5_1, s5_2, s5_3, i4, i5, s4_1, s4_2, s4_3);
s5 : cf_fft_4096_18_5 port map (clock_c, s6_1, s6_2, s6_3, i4, i5, s5_1, s5_2, s5_3);
s6 : cf_fft_4096_18_2 port map (clock_c, i1, i2, i3, i4, i5, s6_1, s6_2, s6_3);
o3 <= s2_3;
o2 <= s2_2;
o1 <= s2_1;
end architecture rtl;

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
entity cf_fft_4096_18 is
port(
signal clock_c : in std_logic;
signal enable_i : in unsigned(0 downto 0);
signal reset_i : in unsigned(0 downto 0);
signal sync_i : in unsigned(0 downto 0);
signal data_0_i : in unsigned(35 downto 0);
signal data_1_i : in unsigned(35 downto 0);
signal sync_o : out unsigned(0 downto 0);
signal data_0_o : out unsigned(35 downto 0);
signal data_1_o : out unsigned(35 downto 0));
end entity cf_fft_4096_18;
architecture rtl of cf_fft_4096_18 is
component cf_fft_4096_18_1 is
port (
clock_c : in std_logic;
i1 : in  unsigned(0 downto 0);
i2 : in  unsigned(35 downto 0);
i3 : in  unsigned(35 downto 0);
i4 : in  unsigned(0 downto 0);
i5 : in  unsigned(0 downto 0);
o1 : out unsigned(0 downto 0);
o2 : out unsigned(35 downto 0);
o3 : out unsigned(35 downto 0));
end component cf_fft_4096_18_1;
signal n1 : unsigned(0 downto 0);
signal n2 : unsigned(35 downto 0);
signal n3 : unsigned(35 downto 0);
begin
s1 : cf_fft_4096_18_1 port map (clock_c, sync_i, data_0_i, data_1_i, enable_i, reset_i, n1, n2, n3);
sync_o <= n1;
data_0_o <= n2;
data_1_o <= n3;
end architecture rtl;


