--
--  Copyright (c) 2003 Launchbird Design Systems, Inc.
--  All rights reserved.
--  
--  Redistribution and use in source and binary forms, with or without modification, are permitted provided that the following conditions are met:
--    Redistributions of source code must retain the above copyright notice, this list of conditions and the following disclaimer.
--    Redistributions in binary form must reproduce the above copyright notice, this list of conditions and the following disclaimer in the documentation and/or other materials provided with the distribution.
--  
--  THIS SOFTWARE IS PROVIDED BY THE COPYRIGHT HOLDERS AND CONTRIBUTORS "AS IS" AND ANY EXPRESS OR IMPLIED WARRANTIES,
--  INCLUDING, BUT NOT LIMITED TO, THE IMPLIED WARRANTIES OF MERCHANTABILITY AND FITNESS FOR A PARTICULAR PURPOSE ARE DISCLAIMED.
--  IN NO EVENT SHALL THE COPYRIGHT OWNER OR CONTRIBUTORS BE LIABLE FOR ANY DIRECT, INDIRECT, INCIDENTAL, SPECIAL, EXEMPLARY,
--  OR CONSEQUENTIAL DAMAGES (INCLUDING, BUT NOT LIMITED TO, PROCUREMENT OF SUBSTITUTE GOODS OR SERVICES; LOSS OF USE, DATA, OR PROFITS;
--  OR BUSINESS INTERRUPTION) HOWEVER CAUSED AND ON ANY THEORY OF LIABILITY, WHETHER IN CONTRACT, STRICT LIABILITY, OR TORT
--  (INCLUDING NEGLIGENCE OR OTHERWISE) ARISING IN ANY WAY OUT OF THE USE OF THIS SOFTWARE, EVEN IF ADVISED OF THE POSSIBILITY OF SUCH DAMAGE.
--  
--  
--  Overview:
--  
--    Performs a radix 2 Fast Fourier Transform.
--    The FFT architecture is pipelined on a rank basis; each rank has its own butterfly and ranks are
--    isolated from each other using memory interleavers.  This FFT can perform calcualations on continuous
--    streaming data (one data set right after another).  More over, inputs and outputs are passed in pairs,
--    doubling the bandwidth.  For instance, a 2048 point FFT can perform a transform every 1024 cycles.
--  
--  Interface:
--  
--    Synchronization:
--      clock_c  : Clock input.
--      enable_i : Synchronous enable.
--      reset_i  : Synchronous reset.
--  
--    Inputs:
--      sync_i     : Input sync pulse must occur one frame prior to data input.
--      data_0_i   : Input data 0.  Width is 2 * precision.  Real on the left, imag on the right.
--      data_1_i   : Input data 1.  Width is 2 * precision.  Real on the left, imag on the right.
--  
--    Outputs:
--      sync_o     : Output sync pulse occurs one frame before data output.
--      data_0_o   : Output data 0.  Width is 2 * precision.  Real on the left, imag on the right.
--      data_1_o   : Output data 1.  Width is 2 * precision.  Real on the left, imag on the right.
--  
--  Built In Parameters:
--  
--    FFT Points   = 256
--    Precision    = 18
--  
--  
--  
--  
--  Generated by Confluence 0.6.3  --  Launchbird Design Systems, Inc.  --  www.launchbird.com
--  
--  Build Date : Fri Aug 22 08:48:47 CDT 2003
--  
--  Interface
--  
--    Build Name    : cf_fft_256_18
--    Clock Domains : clock_c  
--    Vector Input  : enable_i(1)
--    Vector Input  : reset_i(1)
--    Vector Input  : sync_i(1)
--    Vector Input  : data_0_i(36)
--    Vector Input  : data_1_i(36)
--    Vector Output : sync_o(1)
--    Vector Output : data_0_o(36)
--    Vector Output : data_1_o(36)
--  
--  
--  

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
entity cf_fft_256_18_35 is
port (
i1 : in  unsigned(0 downto 0);
i2 : in  unsigned(0 downto 0);
i3 : in  unsigned(0 downto 0);
i4 : in  unsigned(0 downto 0);
i5 : in  unsigned(2 downto 0);
o1 : out unsigned(0 downto 0));
end entity cf_fft_256_18_35;
architecture rtl of cf_fft_256_18_35 is
signal n1 : unsigned(2 downto 0);
signal n2 : unsigned(2 downto 0);
signal n3 : unsigned(2 downto 0);
signal n4 : unsigned(0 downto 0);
signal n5 : unsigned(0 downto 0);
signal n6 : unsigned(0 downto 0);
signal n7 : unsigned(0 downto 0);
signal n8 : unsigned(0 downto 0);
signal n9 : unsigned(0 downto 0);
begin
n1 <= "001";
n2 <= "011";
n3 <= "101";
n4 <= "1" when i5 = n1 else "0";
n5 <= "1" when i5 = n2 else "0";
n6 <= "1" when i5 = n3 else "0";
n7 <= i2 when n6 = "1" else i1;
n8 <= i3 when n5 = "1" else n7;
n9 <= i4 when n4 = "1" else n8;
o1 <= n9;
end architecture rtl;

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
entity cf_fft_256_18_34 is
port (
i1 : in  unsigned(0 downto 0);
i2 : in  unsigned(0 downto 0);
i3 : in  unsigned(0 downto 0);
i4 : in  unsigned(0 downto 0);
i5 : in  unsigned(0 downto 0);
i6 : in  unsigned(0 downto 0);
i7 : in  unsigned(0 downto 0);
i8 : in  unsigned(2 downto 0);
o1 : out unsigned(0 downto 0));
end entity cf_fft_256_18_34;
architecture rtl of cf_fft_256_18_34 is
signal n1 : unsigned(2 downto 0);
signal n2 : unsigned(2 downto 0);
signal n3 : unsigned(2 downto 0);
signal n4 : unsigned(0 downto 0);
signal n5 : unsigned(0 downto 0);
signal n6 : unsigned(0 downto 0);
signal n7 : unsigned(0 downto 0);
signal n8 : unsigned(0 downto 0);
signal n9 : unsigned(0 downto 0);
signal s10_1 : unsigned(0 downto 0);
component cf_fft_256_18_35 is
port (
i1 : in  unsigned(0 downto 0);
i2 : in  unsigned(0 downto 0);
i3 : in  unsigned(0 downto 0);
i4 : in  unsigned(0 downto 0);
i5 : in  unsigned(2 downto 0);
o1 : out unsigned(0 downto 0));
end component cf_fft_256_18_35;
begin
n1 <= "010";
n2 <= "100";
n3 <= "110";
n4 <= "1" when i8 = n1 else "0";
n5 <= "1" when i8 = n2 else "0";
n6 <= "1" when i8 = n3 else "0";
n7 <= i5 when n6 = "1" else s10_1;
n8 <= i6 when n5 = "1" else n7;
n9 <= i7 when n4 = "1" else n8;
s10 : cf_fft_256_18_35 port map (i1, i2, i3, i4, i8, s10_1);
o1 <= n9;
end architecture rtl;

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
entity cf_fft_256_18_33 is
port (
o1 : out unsigned(0 downto 0);
o2 : out unsigned(0 downto 0);
o3 : out unsigned(0 downto 0);
o4 : out unsigned(0 downto 0);
o5 : out unsigned(0 downto 0);
o6 : out unsigned(0 downto 0);
o7 : out unsigned(0 downto 0);
o8 : out unsigned(0 downto 0));
end entity cf_fft_256_18_33;
architecture rtl of cf_fft_256_18_33 is
signal n1 : unsigned(0 downto 0);
signal n2 : unsigned(0 downto 0);
signal n3 : unsigned(0 downto 0);
signal n4 : unsigned(0 downto 0);
signal n5 : unsigned(0 downto 0);
signal n6 : unsigned(0 downto 0);
signal n7 : unsigned(0 downto 0);
signal n8 : unsigned(0 downto 0);
begin
n1 <= "0";
n2 <= "1";
n3 <= "0";
n4 <= "1";
n5 <= "0";
n6 <= "1";
n7 <= "0";
n8 <= "0";
o8 <= n8;
o7 <= n7;
o6 <= n6;
o5 <= n5;
o4 <= n4;
o3 <= n3;
o2 <= n2;
o1 <= n1;
end architecture rtl;

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
entity cf_fft_256_18_32 is
port (
i1 : in  unsigned(0 downto 0);
i2 : in  unsigned(0 downto 0);
i3 : in  unsigned(0 downto 0);
i4 : in  unsigned(2 downto 0);
o1 : out unsigned(0 downto 0));
end entity cf_fft_256_18_32;
architecture rtl of cf_fft_256_18_32 is
signal n1 : unsigned(2 downto 0);
signal n2 : unsigned(2 downto 0);
signal n3 : unsigned(2 downto 0);
signal n4 : unsigned(0 downto 0);
signal n5 : unsigned(0 downto 0);
signal n6 : unsigned(0 downto 0);
signal n7 : unsigned(0 downto 0);
signal n8 : unsigned(0 downto 0);
signal n9 : unsigned(0 downto 0);
signal n10 : unsigned(0 downto 0);
begin
n1 <= "010";
n2 <= "100";
n3 <= "110";
n4 <= "1" when i4 = n1 else "0";
n5 <= "1" when i4 = n2 else "0";
n6 <= "1" when i4 = n3 else "0";
n7 <= i1 when n6 = "1" else n10;
n8 <= i2 when n5 = "1" else n7;
n9 <= i3 when n4 = "1" else n8;
n10 <= "1";
o1 <= n9;
end architecture rtl;

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
entity cf_fft_256_18_31 is
port (
i1 : in  unsigned(2 downto 0);
o1 : out unsigned(0 downto 0));
end entity cf_fft_256_18_31;
architecture rtl of cf_fft_256_18_31 is
signal n1 : unsigned(0 downto 0);
signal n2 : unsigned(0 downto 0);
signal n3 : unsigned(0 downto 0);
signal n4 : unsigned(0 downto 0);
signal n5 : unsigned(2 downto 0);
signal n6 : unsigned(0 downto 0);
signal n7 : unsigned(0 downto 0);
signal s8_1 : unsigned(0 downto 0);
component cf_fft_256_18_32 is
port (
i1 : in  unsigned(0 downto 0);
i2 : in  unsigned(0 downto 0);
i3 : in  unsigned(0 downto 0);
i4 : in  unsigned(2 downto 0);
o1 : out unsigned(0 downto 0));
end component cf_fft_256_18_32;
begin
n1 <= "0";
n2 <= "0";
n3 <= "0";
n4 <= "0";
n5 <= "000";
n6 <= "1" when i1 = n5 else "0";
n7 <= n4 when n6 = "1" else s8_1;
s8 : cf_fft_256_18_32 port map (n1, n2, n3, i1, s8_1);
o1 <= n7;
end architecture rtl;

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
entity cf_fft_256_18_30 is
port (
clock_c : in std_logic;
i1 : in  unsigned(1 downto 0);
i2 : in  unsigned(0 downto 0);
i3 : in  unsigned(0 downto 0);
o1 : out unsigned(0 downto 0));
end entity cf_fft_256_18_30;
architecture rtl of cf_fft_256_18_30 is
signal n1 : unsigned(2 downto 0);
signal n2 : unsigned(2 downto 0);
signal n3 : unsigned(0 downto 0);
signal n4 : unsigned(0 downto 0);
signal n5 : unsigned(0 downto 0) := "0";
signal s6_1 : unsigned(0 downto 0);
signal s7_1 : unsigned(0 downto 0);
signal s7_2 : unsigned(0 downto 0);
signal s7_3 : unsigned(0 downto 0);
signal s7_4 : unsigned(0 downto 0);
signal s7_5 : unsigned(0 downto 0);
signal s7_6 : unsigned(0 downto 0);
signal s7_7 : unsigned(0 downto 0);
signal s7_8 : unsigned(0 downto 0);
signal s8_1 : unsigned(0 downto 0);
component cf_fft_256_18_34 is
port (
i1 : in  unsigned(0 downto 0);
i2 : in  unsigned(0 downto 0);
i3 : in  unsigned(0 downto 0);
i4 : in  unsigned(0 downto 0);
i5 : in  unsigned(0 downto 0);
i6 : in  unsigned(0 downto 0);
i7 : in  unsigned(0 downto 0);
i8 : in  unsigned(2 downto 0);
o1 : out unsigned(0 downto 0));
end component cf_fft_256_18_34;
component cf_fft_256_18_33 is
port (
o1 : out unsigned(0 downto 0);
o2 : out unsigned(0 downto 0);
o3 : out unsigned(0 downto 0);
o4 : out unsigned(0 downto 0);
o5 : out unsigned(0 downto 0);
o6 : out unsigned(0 downto 0);
o7 : out unsigned(0 downto 0);
o8 : out unsigned(0 downto 0));
end component cf_fft_256_18_33;
component cf_fft_256_18_31 is
port (
i1 : in  unsigned(2 downto 0);
o1 : out unsigned(0 downto 0));
end component cf_fft_256_18_31;
begin
n1 <= "000";
n2 <= i1 & n5;
n3 <= "1" when n2 = n1 else "0";
n4 <= s7_8 when n3 = "1" else s6_1;
process (clock_c) begin
  if rising_edge(clock_c) then
    if i3 = "1" then
      n5 <= "0";
    elsif i2 = "1" then
      n5 <= n4;
    end if;
  end if;
end process;
s6 : cf_fft_256_18_34 port map (s7_1, s7_2, s7_3, s7_4, s7_5, s7_6, s7_7, n2, s6_1);
s7 : cf_fft_256_18_33 port map (s7_1, s7_2, s7_3, s7_4, s7_5, s7_6, s7_7, s7_8);
s8 : cf_fft_256_18_31 port map (n2, s8_1);
o1 <= s8_1;
end architecture rtl;

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
entity cf_fft_256_18_29 is
port (
i1 : in  unsigned(0 downto 0);
i2 : in  unsigned(0 downto 0);
i3 : in  unsigned(0 downto 0);
i4 : in  unsigned(0 downto 0);
i5 : in  unsigned(1 downto 0);
o1 : out unsigned(0 downto 0));
end entity cf_fft_256_18_29;
architecture rtl of cf_fft_256_18_29 is
signal n1 : unsigned(1 downto 0);
signal n2 : unsigned(1 downto 0);
signal n3 : unsigned(1 downto 0);
signal n4 : unsigned(0 downto 0);
signal n5 : unsigned(0 downto 0);
signal n6 : unsigned(0 downto 0);
signal n7 : unsigned(0 downto 0);
signal n8 : unsigned(0 downto 0);
signal n9 : unsigned(0 downto 0);
begin
n1 <= "00";
n2 <= "10";
n3 <= "01";
n4 <= "1" when i5 = n1 else "0";
n5 <= "1" when i5 = n2 else "0";
n6 <= "1" when i5 = n3 else "0";
n7 <= i2 when n6 = "1" else i1;
n8 <= i3 when n5 = "1" else n7;
n9 <= i4 when n4 = "1" else n8;
o1 <= n9;
end architecture rtl;

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
entity cf_fft_256_18_28 is
port (
i1 : in  unsigned(1 downto 0);
o1 : out unsigned(0 downto 0));
end entity cf_fft_256_18_28;
architecture rtl of cf_fft_256_18_28 is
signal n1 : unsigned(0 downto 0);
signal n2 : unsigned(0 downto 0);
signal n3 : unsigned(1 downto 0);
signal n4 : unsigned(1 downto 0);
signal n5 : unsigned(0 downto 0);
signal n6 : unsigned(0 downto 0);
signal n7 : unsigned(0 downto 0);
signal n8 : unsigned(0 downto 0);
signal n9 : unsigned(0 downto 0);
begin
n1 <= "0";
n2 <= "0";
n3 <= "00";
n4 <= "10";
n5 <= "1" when i1 = n3 else "0";
n6 <= "1" when i1 = n4 else "0";
n7 <= n1 when n6 = "1" else n9;
n8 <= n2 when n5 = "1" else n7;
n9 <= "1";
o1 <= n8;
end architecture rtl;

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
entity cf_fft_256_18_27 is
port (
clock_c : in std_logic;
i1 : in  unsigned(0 downto 0);
i2 : in  unsigned(0 downto 0);
i3 : in  unsigned(0 downto 0);
o1 : out unsigned(0 downto 0));
end entity cf_fft_256_18_27;
architecture rtl of cf_fft_256_18_27 is
signal n1 : unsigned(0 downto 0);
signal n2 : unsigned(0 downto 0);
signal n3 : unsigned(0 downto 0);
signal n4 : unsigned(0 downto 0);
signal n5 : unsigned(1 downto 0);
signal n6 : unsigned(0 downto 0) := "0";
signal s7_1 : unsigned(0 downto 0);
signal s8_1 : unsigned(0 downto 0);
component cf_fft_256_18_29 is
port (
i1 : in  unsigned(0 downto 0);
i2 : in  unsigned(0 downto 0);
i3 : in  unsigned(0 downto 0);
i4 : in  unsigned(0 downto 0);
i5 : in  unsigned(1 downto 0);
o1 : out unsigned(0 downto 0));
end component cf_fft_256_18_29;
component cf_fft_256_18_28 is
port (
i1 : in  unsigned(1 downto 0);
o1 : out unsigned(0 downto 0));
end component cf_fft_256_18_28;
begin
n1 <= "0";
n2 <= "1";
n3 <= "1";
n4 <= "0";
n5 <= i1 & n6;
process (clock_c) begin
  if rising_edge(clock_c) then
    if i3 = "1" then
      n6 <= "0";
    elsif i2 = "1" then
      n6 <= s7_1;
    end if;
  end if;
end process;
s7 : cf_fft_256_18_29 port map (n1, n2, n3, n4, n5, s7_1);
s8 : cf_fft_256_18_28 port map (n5, s8_1);
o1 <= s8_1;
end architecture rtl;

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
entity cf_fft_256_18_26 is
port (
clock_c : in std_logic;
i1 : in  unsigned(0 downto 0);
i2 : in  unsigned(71 downto 0);
i3 : in  unsigned(0 downto 0);
i4 : in  unsigned(5 downto 0);
i5 : in  unsigned(0 downto 0);
i6 : in  unsigned(0 downto 0);
o1 : out unsigned(71 downto 0));
end entity cf_fft_256_18_26;
architecture rtl of cf_fft_256_18_26 is
signal n1 : unsigned(5 downto 0);
signal n2 : unsigned(5 downto 0);
signal n3 : unsigned(5 downto 0) := "000000";
signal n4 : unsigned(0 downto 0);
signal n5 : unsigned(0 downto 0);
signal n6 : unsigned(71 downto 0);
signal n6a : unsigned(5 downto 0) := "000000";
type   n6mt is array (63 downto 0) of unsigned(71 downto 0);
signal n6m : n6mt;
signal n7 : unsigned(0 downto 0);
signal n8 : unsigned(71 downto 0);
signal n8a : unsigned(5 downto 0) := "000000";
type   n8mt is array (63 downto 0) of unsigned(71 downto 0);
signal n8m : n8mt;
signal n9 : unsigned(0 downto 0) := "0";
signal n10 : unsigned(71 downto 0);
signal n11 : unsigned(0 downto 0);
signal s12_1 : unsigned(0 downto 0);
component cf_fft_256_18_27 is
port (
clock_c : in std_logic;
i1 : in  unsigned(0 downto 0);
i2 : in  unsigned(0 downto 0);
i3 : in  unsigned(0 downto 0);
o1 : out unsigned(0 downto 0));
end component cf_fft_256_18_27;
begin
n1 <= "000001";
n2 <= n3 + n1;
process (clock_c) begin
  if rising_edge(clock_c) then
    if n11 = "1" then
      n3 <= "000000";
    elsif i5 = "1" then
      n3 <= n2;
    end if;
  end if;
end process;
n4 <= not s12_1;
n5 <= i3 and n4;
process (clock_c) begin
  if rising_edge(clock_c) then
    if i5 = "1" then
      if n5 = "1" then
        n6m(to_integer(i4)) <= i2;
      end if;
      n6a <= n3;
    end if;
  end if;
end process;
n6 <= n6m(to_integer(n6a));
n7 <= i3 and s12_1;
process (clock_c) begin
  if rising_edge(clock_c) then
    if i5 = "1" then
      if n7 = "1" then
        n8m(to_integer(i4)) <= i2;
      end if;
      n8a <= n3;
    end if;
  end if;
end process;
n8 <= n8m(to_integer(n8a));
process (clock_c) begin
  if rising_edge(clock_c) then
    if i6 = "1" then
      n9 <= "0";
    elsif i5 = "1" then
      n9 <= n4;
    end if;
  end if;
end process;
n10 <= n8 when n9 = "1" else n6;
n11 <= i1 or i6;
s12 : cf_fft_256_18_27 port map (clock_c, i1, i5, i6, s12_1);
o1 <= n10;
end architecture rtl;

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
entity cf_fft_256_18_25 is
port (
clock_c : in std_logic;
i1 : in  unsigned(0 downto 0);
i2 : in  unsigned(71 downto 0);
i3 : in  unsigned(0 downto 0);
i4 : in  unsigned(5 downto 0);
i5 : in  unsigned(0 downto 0);
i6 : in  unsigned(0 downto 0);
o1 : out unsigned(0 downto 0);
o2 : out unsigned(0 downto 0);
o3 : out unsigned(71 downto 0));
end entity cf_fft_256_18_25;
architecture rtl of cf_fft_256_18_25 is
signal n1 : unsigned(5 downto 0);
signal n2 : unsigned(5 downto 0);
signal n3 : unsigned(5 downto 0) := "000000";
signal n4 : unsigned(0 downto 0);
signal n5 : unsigned(0 downto 0) := "0";
signal n6 : unsigned(5 downto 0);
signal n7 : unsigned(0 downto 0);
signal n8 : unsigned(0 downto 0);
signal n9 : unsigned(71 downto 0);
signal n9a : unsigned(5 downto 0) := "000000";
type   n9mt is array (63 downto 0) of unsigned(71 downto 0);
signal n9m : n9mt;
signal n10 : unsigned(0 downto 0);
signal n11 : unsigned(71 downto 0);
signal n11a : unsigned(5 downto 0) := "000000";
type   n11mt is array (63 downto 0) of unsigned(71 downto 0);
signal n11m : n11mt;
signal n12 : unsigned(0 downto 0) := "0";
signal n13 : unsigned(71 downto 0);
signal n14 : unsigned(0 downto 0);
signal s15_1 : unsigned(0 downto 0);
component cf_fft_256_18_27 is
port (
clock_c : in std_logic;
i1 : in  unsigned(0 downto 0);
i2 : in  unsigned(0 downto 0);
i3 : in  unsigned(0 downto 0);
o1 : out unsigned(0 downto 0));
end component cf_fft_256_18_27;
begin
n1 <= "000001";
n2 <= n3 + n1;
process (clock_c) begin
  if rising_edge(clock_c) then
    if n14 = "1" then
      n3 <= "000000";
    elsif i5 = "1" then
      n3 <= n2;
    end if;
  end if;
end process;
n4 <= not s15_1;
process (clock_c) begin
  if rising_edge(clock_c) then
    if i6 = "1" then
      n5 <= "0";
    elsif i5 = "1" then
      n5 <= i1;
    end if;
  end if;
end process;
n6 <= "000000";
n7 <= "1" when n3 = n6 else "0";
n8 <= i3 and n4;
process (clock_c) begin
  if rising_edge(clock_c) then
    if i5 = "1" then
      if n8 = "1" then
        n9m(to_integer(i4)) <= i2;
      end if;
      n9a <= n3;
    end if;
  end if;
end process;
n9 <= n9m(to_integer(n9a));
n10 <= i3 and s15_1;
process (clock_c) begin
  if rising_edge(clock_c) then
    if i5 = "1" then
      if n10 = "1" then
        n11m(to_integer(i4)) <= i2;
      end if;
      n11a <= n3;
    end if;
  end if;
end process;
n11 <= n11m(to_integer(n11a));
process (clock_c) begin
  if rising_edge(clock_c) then
    if i6 = "1" then
      n12 <= "0";
    elsif i5 = "1" then
      n12 <= n4;
    end if;
  end if;
end process;
n13 <= n11 when n12 = "1" else n9;
n14 <= i1 or i6;
s15 : cf_fft_256_18_27 port map (clock_c, i1, i5, i6, s15_1);
o3 <= n13;
o2 <= n7;
o1 <= n5;
end architecture rtl;

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
entity cf_fft_256_18_24 is
port (
i1 : in  unsigned(0 downto 0);
i2 : in  unsigned(0 downto 0);
i3 : in  unsigned(0 downto 0);
i4 : in  unsigned(2 downto 0);
o1 : out unsigned(0 downto 0));
end entity cf_fft_256_18_24;
architecture rtl of cf_fft_256_18_24 is
signal n1 : unsigned(2 downto 0);
signal n2 : unsigned(2 downto 0);
signal n3 : unsigned(2 downto 0);
signal n4 : unsigned(0 downto 0);
signal n5 : unsigned(0 downto 0);
signal n6 : unsigned(0 downto 0);
signal n7 : unsigned(0 downto 0);
signal n8 : unsigned(0 downto 0);
signal n9 : unsigned(0 downto 0);
signal n10 : unsigned(0 downto 0);
begin
n1 <= "110";
n2 <= "001";
n3 <= "011";
n4 <= "1" when i4 = n1 else "0";
n5 <= "1" when i4 = n2 else "0";
n6 <= "1" when i4 = n3 else "0";
n7 <= i1 when n6 = "1" else n10;
n8 <= i2 when n5 = "1" else n7;
n9 <= i3 when n4 = "1" else n8;
n10 <= "1";
o1 <= n9;
end architecture rtl;

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
entity cf_fft_256_18_23 is
port (
i1 : in  unsigned(0 downto 0);
i2 : in  unsigned(0 downto 0);
i3 : in  unsigned(0 downto 0);
i4 : in  unsigned(0 downto 0);
i5 : in  unsigned(0 downto 0);
i6 : in  unsigned(0 downto 0);
i7 : in  unsigned(2 downto 0);
o1 : out unsigned(0 downto 0));
end entity cf_fft_256_18_23;
architecture rtl of cf_fft_256_18_23 is
signal n1 : unsigned(2 downto 0);
signal n2 : unsigned(2 downto 0);
signal n3 : unsigned(2 downto 0);
signal n4 : unsigned(0 downto 0);
signal n5 : unsigned(0 downto 0);
signal n6 : unsigned(0 downto 0);
signal n7 : unsigned(0 downto 0);
signal n8 : unsigned(0 downto 0);
signal n9 : unsigned(0 downto 0);
signal s10_1 : unsigned(0 downto 0);
component cf_fft_256_18_24 is
port (
i1 : in  unsigned(0 downto 0);
i2 : in  unsigned(0 downto 0);
i3 : in  unsigned(0 downto 0);
i4 : in  unsigned(2 downto 0);
o1 : out unsigned(0 downto 0));
end component cf_fft_256_18_24;
begin
n1 <= "000";
n2 <= "010";
n3 <= "100";
n4 <= "1" when i7 = n1 else "0";
n5 <= "1" when i7 = n2 else "0";
n6 <= "1" when i7 = n3 else "0";
n7 <= i4 when n6 = "1" else s10_1;
n8 <= i5 when n5 = "1" else n7;
n9 <= i6 when n4 = "1" else n8;
s10 : cf_fft_256_18_24 port map (i1, i2, i3, i7, s10_1);
o1 <= n9;
end architecture rtl;

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
entity cf_fft_256_18_22 is
port (
clock_c : in std_logic;
i1 : in  unsigned(1 downto 0);
i2 : in  unsigned(0 downto 0);
i3 : in  unsigned(0 downto 0);
o1 : out unsigned(0 downto 0));
end entity cf_fft_256_18_22;
architecture rtl of cf_fft_256_18_22 is
signal n1 : unsigned(0 downto 0);
signal n2 : unsigned(0 downto 0);
signal n3 : unsigned(0 downto 0);
signal n4 : unsigned(0 downto 0);
signal n5 : unsigned(0 downto 0);
signal n6 : unsigned(0 downto 0);
signal n7 : unsigned(0 downto 0);
signal n8 : unsigned(0 downto 0);
signal n9 : unsigned(0 downto 0);
signal n10 : unsigned(0 downto 0);
signal n11 : unsigned(0 downto 0);
signal n12 : unsigned(0 downto 0);
signal n13 : unsigned(2 downto 0);
signal n14 : unsigned(0 downto 0) := "0";
signal s15_1 : unsigned(0 downto 0);
signal s16_1 : unsigned(0 downto 0);
component cf_fft_256_18_23 is
port (
i1 : in  unsigned(0 downto 0);
i2 : in  unsigned(0 downto 0);
i3 : in  unsigned(0 downto 0);
i4 : in  unsigned(0 downto 0);
i5 : in  unsigned(0 downto 0);
i6 : in  unsigned(0 downto 0);
i7 : in  unsigned(2 downto 0);
o1 : out unsigned(0 downto 0));
end component cf_fft_256_18_23;
begin
n1 <= "0";
n2 <= "1";
n3 <= "1";
n4 <= "1";
n5 <= "0";
n6 <= "0";
n7 <= "0";
n8 <= "1";
n9 <= "1";
n10 <= "1";
n11 <= "0";
n12 <= "0";
n13 <= i1 & n14;
process (clock_c) begin
  if rising_edge(clock_c) then
    if i3 = "1" then
      n14 <= "0";
    elsif i2 = "1" then
      n14 <= s15_1;
    end if;
  end if;
end process;
s15 : cf_fft_256_18_23 port map (n1, n2, n3, n4, n5, n6, n13, s15_1);
s16 : cf_fft_256_18_23 port map (n7, n8, n9, n10, n11, n12, n13, s16_1);
o1 <= s16_1;
end architecture rtl;

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
entity cf_fft_256_18_21 is
port (
clock_c : in std_logic;
i1 : in  unsigned(0 downto 0);
i2 : in  unsigned(0 downto 0);
i3 : in  unsigned(0 downto 0);
o1 : out unsigned(6 downto 0);
o2 : out unsigned(0 downto 0));
end entity cf_fft_256_18_21;
architecture rtl of cf_fft_256_18_21 is
signal n1 : unsigned(6 downto 0);
signal n2 : unsigned(6 downto 0);
signal n3 : unsigned(6 downto 0) := "0000000";
signal n4 : unsigned(6 downto 0);
signal n5 : unsigned(0 downto 0);
signal n6 : unsigned(1 downto 0);
signal n7 : unsigned(0 downto 0) := "0";
signal n8 : unsigned(0 downto 0);
signal n9 : unsigned(0 downto 0);
signal n10 : unsigned(0 downto 0);
signal s11_1 : unsigned(0 downto 0);
component cf_fft_256_18_22 is
port (
clock_c : in std_logic;
i1 : in  unsigned(1 downto 0);
i2 : in  unsigned(0 downto 0);
i3 : in  unsigned(0 downto 0);
o1 : out unsigned(0 downto 0));
end component cf_fft_256_18_22;
begin
n1 <= "0000001";
n2 <= n3 + n1;
process (clock_c) begin
  if rising_edge(clock_c) then
    if n9 = "1" then
      n3 <= "0000000";
    elsif n10 = "1" then
      n3 <= n2;
    end if;
  end if;
end process;
n4 <= "1111111";
n5 <= "1" when n3 = n4 else "0";
n6 <= i1 & n5;
process (clock_c) begin
  if rising_edge(clock_c) then
    if i3 = "1" then
      n7 <= "0";
    elsif i2 = "1" then
      n7 <= s11_1;
    end if;
  end if;
end process;
n8 <= n7 and n5;
n9 <= i1 or i3;
n10 <= s11_1 and i2;
s11 : cf_fft_256_18_22 port map (clock_c, n6, i2, i3, s11_1);
o2 <= n8;
o1 <= n3;
end architecture rtl;

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
entity cf_fft_256_18_20 is
port (
clock_c : in std_logic;
i1 : in  unsigned(0 downto 0);
i2 : in  unsigned(35 downto 0);
i3 : in  unsigned(35 downto 0);
i4 : in  unsigned(0 downto 0);
i5 : in  unsigned(0 downto 0);
o1 : out unsigned(0 downto 0);
o2 : out unsigned(35 downto 0);
o3 : out unsigned(35 downto 0));
end entity cf_fft_256_18_20;
architecture rtl of cf_fft_256_18_20 is
signal n1 : unsigned(71 downto 0);
signal n2 : unsigned(0 downto 0);
signal n3 : unsigned(0 downto 0);
signal n4 : unsigned(5 downto 0);
signal n5 : unsigned(5 downto 0);
signal n6 : unsigned(1 downto 0);
signal n7 : unsigned(35 downto 0);
signal n8 : unsigned(35 downto 0);
signal n9 : unsigned(35 downto 0);
signal n10 : unsigned(35 downto 0);
signal n11 : unsigned(35 downto 0);
signal n12 : unsigned(35 downto 0);
signal s13_1 : unsigned(0 downto 0);
signal s14_1 : unsigned(71 downto 0);
signal s15_1 : unsigned(0 downto 0);
signal s15_2 : unsigned(0 downto 0);
signal s15_3 : unsigned(71 downto 0);
signal s16_1 : unsigned(6 downto 0);
signal s16_2 : unsigned(0 downto 0);
component cf_fft_256_18_30 is
port (
clock_c : in std_logic;
i1 : in  unsigned(1 downto 0);
i2 : in  unsigned(0 downto 0);
i3 : in  unsigned(0 downto 0);
o1 : out unsigned(0 downto 0));
end component cf_fft_256_18_30;
component cf_fft_256_18_26 is
port (
clock_c : in std_logic;
i1 : in  unsigned(0 downto 0);
i2 : in  unsigned(71 downto 0);
i3 : in  unsigned(0 downto 0);
i4 : in  unsigned(5 downto 0);
i5 : in  unsigned(0 downto 0);
i6 : in  unsigned(0 downto 0);
o1 : out unsigned(71 downto 0));
end component cf_fft_256_18_26;
component cf_fft_256_18_25 is
port (
clock_c : in std_logic;
i1 : in  unsigned(0 downto 0);
i2 : in  unsigned(71 downto 0);
i3 : in  unsigned(0 downto 0);
i4 : in  unsigned(5 downto 0);
i5 : in  unsigned(0 downto 0);
i6 : in  unsigned(0 downto 0);
o1 : out unsigned(0 downto 0);
o2 : out unsigned(0 downto 0);
o3 : out unsigned(71 downto 0));
end component cf_fft_256_18_25;
component cf_fft_256_18_21 is
port (
clock_c : in std_logic;
i1 : in  unsigned(0 downto 0);
i2 : in  unsigned(0 downto 0);
i3 : in  unsigned(0 downto 0);
o1 : out unsigned(6 downto 0);
o2 : out unsigned(0 downto 0));
end component cf_fft_256_18_21;
begin
n1 <= i2 & i3;
n2 <= s16_1(6 downto 6);
n3 <= not n2;
n4 <= s16_1(5 downto 5) &
  s16_1(4 downto 4) &
  s16_1(3 downto 3) &
  s16_1(2 downto 2) &
  s16_1(1 downto 1) &
  s16_1(0 downto 0);
n5 <= n4(0 downto 0) &
  n4(1 downto 1) &
  n4(2 downto 2) &
  n4(3 downto 3) &
  n4(4 downto 4) &
  n4(5 downto 5);
n6 <= s15_2 & s15_1;
n7 <= s15_3(71 downto 71) &
  s15_3(70 downto 70) &
  s15_3(69 downto 69) &
  s15_3(68 downto 68) &
  s15_3(67 downto 67) &
  s15_3(66 downto 66) &
  s15_3(65 downto 65) &
  s15_3(64 downto 64) &
  s15_3(63 downto 63) &
  s15_3(62 downto 62) &
  s15_3(61 downto 61) &
  s15_3(60 downto 60) &
  s15_3(59 downto 59) &
  s15_3(58 downto 58) &
  s15_3(57 downto 57) &
  s15_3(56 downto 56) &
  s15_3(55 downto 55) &
  s15_3(54 downto 54) &
  s15_3(53 downto 53) &
  s15_3(52 downto 52) &
  s15_3(51 downto 51) &
  s15_3(50 downto 50) &
  s15_3(49 downto 49) &
  s15_3(48 downto 48) &
  s15_3(47 downto 47) &
  s15_3(46 downto 46) &
  s15_3(45 downto 45) &
  s15_3(44 downto 44) &
  s15_3(43 downto 43) &
  s15_3(42 downto 42) &
  s15_3(41 downto 41) &
  s15_3(40 downto 40) &
  s15_3(39 downto 39) &
  s15_3(38 downto 38) &
  s15_3(37 downto 37) &
  s15_3(36 downto 36);
n8 <= s15_3(35 downto 35) &
  s15_3(34 downto 34) &
  s15_3(33 downto 33) &
  s15_3(32 downto 32) &
  s15_3(31 downto 31) &
  s15_3(30 downto 30) &
  s15_3(29 downto 29) &
  s15_3(28 downto 28) &
  s15_3(27 downto 27) &
  s15_3(26 downto 26) &
  s15_3(25 downto 25) &
  s15_3(24 downto 24) &
  s15_3(23 downto 23) &
  s15_3(22 downto 22) &
  s15_3(21 downto 21) &
  s15_3(20 downto 20) &
  s15_3(19 downto 19) &
  s15_3(18 downto 18) &
  s15_3(17 downto 17) &
  s15_3(16 downto 16) &
  s15_3(15 downto 15) &
  s15_3(14 downto 14) &
  s15_3(13 downto 13) &
  s15_3(12 downto 12) &
  s15_3(11 downto 11) &
  s15_3(10 downto 10) &
  s15_3(9 downto 9) &
  s15_3(8 downto 8) &
  s15_3(7 downto 7) &
  s15_3(6 downto 6) &
  s15_3(5 downto 5) &
  s15_3(4 downto 4) &
  s15_3(3 downto 3) &
  s15_3(2 downto 2) &
  s15_3(1 downto 1) &
  s15_3(0 downto 0);
n9 <= s14_1(71 downto 71) &
  s14_1(70 downto 70) &
  s14_1(69 downto 69) &
  s14_1(68 downto 68) &
  s14_1(67 downto 67) &
  s14_1(66 downto 66) &
  s14_1(65 downto 65) &
  s14_1(64 downto 64) &
  s14_1(63 downto 63) &
  s14_1(62 downto 62) &
  s14_1(61 downto 61) &
  s14_1(60 downto 60) &
  s14_1(59 downto 59) &
  s14_1(58 downto 58) &
  s14_1(57 downto 57) &
  s14_1(56 downto 56) &
  s14_1(55 downto 55) &
  s14_1(54 downto 54) &
  s14_1(53 downto 53) &
  s14_1(52 downto 52) &
  s14_1(51 downto 51) &
  s14_1(50 downto 50) &
  s14_1(49 downto 49) &
  s14_1(48 downto 48) &
  s14_1(47 downto 47) &
  s14_1(46 downto 46) &
  s14_1(45 downto 45) &
  s14_1(44 downto 44) &
  s14_1(43 downto 43) &
  s14_1(42 downto 42) &
  s14_1(41 downto 41) &
  s14_1(40 downto 40) &
  s14_1(39 downto 39) &
  s14_1(38 downto 38) &
  s14_1(37 downto 37) &
  s14_1(36 downto 36);
n10 <= s14_1(35 downto 35) &
  s14_1(34 downto 34) &
  s14_1(33 downto 33) &
  s14_1(32 downto 32) &
  s14_1(31 downto 31) &
  s14_1(30 downto 30) &
  s14_1(29 downto 29) &
  s14_1(28 downto 28) &
  s14_1(27 downto 27) &
  s14_1(26 downto 26) &
  s14_1(25 downto 25) &
  s14_1(24 downto 24) &
  s14_1(23 downto 23) &
  s14_1(22 downto 22) &
  s14_1(21 downto 21) &
  s14_1(20 downto 20) &
  s14_1(19 downto 19) &
  s14_1(18 downto 18) &
  s14_1(17 downto 17) &
  s14_1(16 downto 16) &
  s14_1(15 downto 15) &
  s14_1(14 downto 14) &
  s14_1(13 downto 13) &
  s14_1(12 downto 12) &
  s14_1(11 downto 11) &
  s14_1(10 downto 10) &
  s14_1(9 downto 9) &
  s14_1(8 downto 8) &
  s14_1(7 downto 7) &
  s14_1(6 downto 6) &
  s14_1(5 downto 5) &
  s14_1(4 downto 4) &
  s14_1(3 downto 3) &
  s14_1(2 downto 2) &
  s14_1(1 downto 1) &
  s14_1(0 downto 0);
n11 <= n8 when s13_1 = "1" else n7;
n12 <= n10 when s13_1 = "1" else n9;
s13 : cf_fft_256_18_30 port map (clock_c, n6, i4, i5, s13_1);
s14 : cf_fft_256_18_26 port map (clock_c, s16_2, n1, n2, n5, i4, i5, s14_1);
s15 : cf_fft_256_18_25 port map (clock_c, s16_2, n1, n3, n5, i4, i5, s15_1, s15_2, s15_3);
s16 : cf_fft_256_18_21 port map (clock_c, i1, i4, i5, s16_1, s16_2);
o3 <= n12;
o2 <= n11;
o1 <= s15_1;
end architecture rtl;

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
entity cf_fft_256_18_19 is
port (
clock_c : in std_logic;
i1 : in  unsigned(35 downto 0);
i2 : in  unsigned(35 downto 0);
i3 : in  unsigned(5 downto 0);
i4 : in  unsigned(0 downto 0);
i5 : in  unsigned(0 downto 0);
o1 : out unsigned(35 downto 0);
o2 : out unsigned(35 downto 0));
end entity cf_fft_256_18_19;
architecture rtl of cf_fft_256_18_19 is
signal n1 : unsigned(35 downto 0) := "000000000000000000000000000000000000";
signal n2 : unsigned(17 downto 0);
signal n3 : unsigned(17 downto 0);
signal n4 : unsigned(35 downto 0) := "000000000000000000000000000000000000";
signal n5 : unsigned(17 downto 0);
signal n6 : unsigned(17 downto 0);
signal n7 : unsigned(17 downto 0) := "000000000000000000";
signal n8 : unsigned(17 downto 0) := "000000000000000000";
signal n9 : unsigned(17 downto 0) := "000000000000000000";
signal n10 : unsigned(17 downto 0) := "000000000000000000";
signal n11 : unsigned(35 downto 0) := "000000000000000000000000000000000000";
signal n12 : unsigned(17 downto 0);
signal n13 : unsigned(17 downto 0);
signal n14 : unsigned(35 downto 0);
signal n15 : unsigned(17 downto 0);
signal n16 : unsigned(17 downto 0) := "000000000000000000";
signal n17 : unsigned(35 downto 0);
signal n18 : unsigned(17 downto 0);
signal n19 : unsigned(17 downto 0) := "000000000000000000";
signal n20 : unsigned(17 downto 0);
signal n21 : unsigned(17 downto 0) := "000000000000000000";
signal n22 : unsigned(35 downto 0);
signal n23 : unsigned(17 downto 0);
signal n24 : unsigned(17 downto 0) := "000000000000000000";
signal n25 : unsigned(35 downto 0);
signal n26 : unsigned(17 downto 0);
signal n27 : unsigned(17 downto 0) := "000000000000000000";
signal n28 : unsigned(17 downto 0);
signal n29 : unsigned(17 downto 0) := "000000000000000000";
signal n30 : unsigned(17 downto 0);
signal n31 : unsigned(17 downto 0);
signal n32 : unsigned(35 downto 0);
signal n33 : unsigned(35 downto 0) := "000000000000000000000000000000000000";
signal n34 : unsigned(17 downto 0);
signal n35 : unsigned(17 downto 0);
signal n36 : unsigned(35 downto 0);
signal n37 : unsigned(35 downto 0) := "000000000000000000000000000000000000";
begin
process (clock_c) begin
  if rising_edge(clock_c) then
    if i5 = "1" then
      n1 <= "000000000000000000000000000000000000";
    elsif i4 = "1" then
      n1 <= i1;
    end if;
  end if;
end process;
n2 <= n1(35 downto 35) &
  n1(34 downto 34) &
  n1(33 downto 33) &
  n1(32 downto 32) &
  n1(31 downto 31) &
  n1(30 downto 30) &
  n1(29 downto 29) &
  n1(28 downto 28) &
  n1(27 downto 27) &
  n1(26 downto 26) &
  n1(25 downto 25) &
  n1(24 downto 24) &
  n1(23 downto 23) &
  n1(22 downto 22) &
  n1(21 downto 21) &
  n1(20 downto 20) &
  n1(19 downto 19) &
  n1(18 downto 18);
n3 <= n1(17 downto 17) &
  n1(16 downto 16) &
  n1(15 downto 15) &
  n1(14 downto 14) &
  n1(13 downto 13) &
  n1(12 downto 12) &
  n1(11 downto 11) &
  n1(10 downto 10) &
  n1(9 downto 9) &
  n1(8 downto 8) &
  n1(7 downto 7) &
  n1(6 downto 6) &
  n1(5 downto 5) &
  n1(4 downto 4) &
  n1(3 downto 3) &
  n1(2 downto 2) &
  n1(1 downto 1) &
  n1(0 downto 0);
process (clock_c) begin
  if rising_edge(clock_c) then
    if i5 = "1" then
      n4 <= "000000000000000000000000000000000000";
    elsif i4 = "1" then
      n4 <= i2;
    end if;
  end if;
end process;
n5 <= n4(35 downto 35) &
  n4(34 downto 34) &
  n4(33 downto 33) &
  n4(32 downto 32) &
  n4(31 downto 31) &
  n4(30 downto 30) &
  n4(29 downto 29) &
  n4(28 downto 28) &
  n4(27 downto 27) &
  n4(26 downto 26) &
  n4(25 downto 25) &
  n4(24 downto 24) &
  n4(23 downto 23) &
  n4(22 downto 22) &
  n4(21 downto 21) &
  n4(20 downto 20) &
  n4(19 downto 19) &
  n4(18 downto 18);
n6 <= n4(17 downto 17) &
  n4(16 downto 16) &
  n4(15 downto 15) &
  n4(14 downto 14) &
  n4(13 downto 13) &
  n4(12 downto 12) &
  n4(11 downto 11) &
  n4(10 downto 10) &
  n4(9 downto 9) &
  n4(8 downto 8) &
  n4(7 downto 7) &
  n4(6 downto 6) &
  n4(5 downto 5) &
  n4(4 downto 4) &
  n4(3 downto 3) &
  n4(2 downto 2) &
  n4(1 downto 1) &
  n4(0 downto 0);
process (clock_c) begin
  if rising_edge(clock_c) then
    if i5 = "1" then
      n7 <= "000000000000000000";
    elsif i4 = "1" then
      n7 <= n2;
    end if;
  end if;
end process;
process (clock_c) begin
  if rising_edge(clock_c) then
    if i5 = "1" then
      n8 <= "000000000000000000";
    elsif i4 = "1" then
      n8 <= n7;
    end if;
  end if;
end process;
process (clock_c) begin
  if rising_edge(clock_c) then
    if i5 = "1" then
      n9 <= "000000000000000000";
    elsif i4 = "1" then
      n9 <= n3;
    end if;
  end if;
end process;
process (clock_c) begin
  if rising_edge(clock_c) then
    if i5 = "1" then
      n10 <= "000000000000000000";
    elsif i4 = "1" then
      n10 <= n9;
    end if;
  end if;
end process;
process (clock_c) begin
  if rising_edge(clock_c) then 
    if i4 = "1" then
      case i3 is
        when "000000" => n11 <= "011111111111111111000000000000000000";
        when "000001" => n11 <= "011111111101100010111110011011100000";
        when "000010" => n11 <= "011111110110001000111100110111010000";
        when "000011" => n11 <= "011111101001110101111011010011011111";
        when "000100" => n11 <= "011111011000101001111001110000011101";
        when "000101" => n11 <= "011111000010100111111000001110011000";
        when "000110" => n11 <= "011110100111110100110110101101011111";
        when "000111" => n11 <= "011110001000010010110101001110000011";
        when "001000" => n11 <= "011101100100000110110011110000010000";
        when "001001" => n11 <= "011100111011010111110010010100010111";
        when "001010" => n11 <= "011100001110001011110000111010100101";
        when "001011" => n11 <= "011011011100101000101111100011000111";
        when "001100" => n11 <= "011010100110110110101110001110001100";
        when "001101" => n11 <= "011001101100111110101100111100000000";
        when "001110" => n11 <= "011000101111001000101011101100110000";
        when "001111" => n11 <= "010111101101011101101010100000101001";
        when "010000" => n11 <= "010110101000001001101001010111110110";
        when "010001" => n11 <= "010101011111010110101000010010100010";
        when "010010" => n11 <= "010100010011001111100111010000110111";
        when "010011" => n11 <= "010011000011111111100110010011000001";
        when "010100" => n11 <= "010001110001110011100101011001001001";
        when "010101" => n11 <= "010000011100111000100100100011010111";
        when "010110" => n11 <= "001111000101011010100011110001110100";
        when "010111" => n11 <= "001101101011101000100011000100101000";
        when "011000" => n11 <= "001100001111101111100010011011111001";
        when "011001" => n11 <= "001010110001111100100001110111101101";
        when "011010" => n11 <= "001001010010100000100001011000001011";
        when "011011" => n11 <= "000111110001100111100000111101011000";
        when "011100" => n11 <= "000110001111100010100000100111010110";
        when "011101" => n11 <= "000100101100100000100000010110001010";
        when "011110" => n11 <= "000011001000101111100000001001110111";
        when "011111" => n11 <= "000001100100011111100000000010011101";
        when "100000" => n11 <= "000000000000000000100000000000000000";
        when "100001" => n11 <= "111110011011100000100000000010011101";
        when "100010" => n11 <= "111100110111010000100000001001110111";
        when "100011" => n11 <= "111011010011011111100000010110001010";
        when "100100" => n11 <= "111001110000011101100000100111010110";
        when "100101" => n11 <= "111000001110011000100000111101011000";
        when "100110" => n11 <= "110110101101011111100001011000001011";
        when "100111" => n11 <= "110101001110000011100001110111101101";
        when "101000" => n11 <= "110011110000010000100010011011111001";
        when "101001" => n11 <= "110010010100010111100011000100101000";
        when "101010" => n11 <= "110000111010100101100011110001110100";
        when "101011" => n11 <= "101111100011000111100100100011010111";
        when "101100" => n11 <= "101110001110001100100101011001001001";
        when "101101" => n11 <= "101100111100000000100110010011000001";
        when "101110" => n11 <= "101011101100110000100111010000110111";
        when "101111" => n11 <= "101010100000101001101000010010100010";
        when "110000" => n11 <= "101001010111110110101001010111110110";
        when "110001" => n11 <= "101000010010100010101010100000101001";
        when "110010" => n11 <= "100111010000110111101011101100110000";
        when "110011" => n11 <= "100110010011000001101100111100000000";
        when "110100" => n11 <= "100101011001001001101110001110001100";
        when "110101" => n11 <= "100100100011010111101111100011000111";
        when "110110" => n11 <= "100011110001110100110000111010100101";
        when "110111" => n11 <= "100011000100101000110010010100010111";
        when "111000" => n11 <= "100010011011111001110011110000010000";
        when "111001" => n11 <= "100001110111101101110101001110000011";
        when "111010" => n11 <= "100001011000001011110110101101011111";
        when "111011" => n11 <= "100000111101011000111000001110011000";
        when "111100" => n11 <= "100000100111010110111001110000011101";
        when "111101" => n11 <= "100000010110001010111011010011011111";
        when "111110" => n11 <= "100000001001110111111100110111010000";
        when "111111" => n11 <= "100000000010011101111110011011100000";
        when others => n11 <= "XXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX";
      end case;
    end if;
  end if;
end process;
n12 <= n11(35 downto 35) &
  n11(34 downto 34) &
  n11(33 downto 33) &
  n11(32 downto 32) &
  n11(31 downto 31) &
  n11(30 downto 30) &
  n11(29 downto 29) &
  n11(28 downto 28) &
  n11(27 downto 27) &
  n11(26 downto 26) &
  n11(25 downto 25) &
  n11(24 downto 24) &
  n11(23 downto 23) &
  n11(22 downto 22) &
  n11(21 downto 21) &
  n11(20 downto 20) &
  n11(19 downto 19) &
  n11(18 downto 18);
n13 <= n11(17 downto 17) &
  n11(16 downto 16) &
  n11(15 downto 15) &
  n11(14 downto 14) &
  n11(13 downto 13) &
  n11(12 downto 12) &
  n11(11 downto 11) &
  n11(10 downto 10) &
  n11(9 downto 9) &
  n11(8 downto 8) &
  n11(7 downto 7) &
  n11(6 downto 6) &
  n11(5 downto 5) &
  n11(4 downto 4) &
  n11(3 downto 3) &
  n11(2 downto 2) &
  n11(1 downto 1) &
  n11(0 downto 0);
n14 <= unsigned(signed(n5) * signed(n12));
n15 <= n14(34 downto 34) &
  n14(33 downto 33) &
  n14(32 downto 32) &
  n14(31 downto 31) &
  n14(30 downto 30) &
  n14(29 downto 29) &
  n14(28 downto 28) &
  n14(27 downto 27) &
  n14(26 downto 26) &
  n14(25 downto 25) &
  n14(24 downto 24) &
  n14(23 downto 23) &
  n14(22 downto 22) &
  n14(21 downto 21) &
  n14(20 downto 20) &
  n14(19 downto 19) &
  n14(18 downto 18) &
  n14(17 downto 17);
process (clock_c) begin
  if rising_edge(clock_c) then
    if i5 = "1" then
      n16 <= "000000000000000000";
    elsif i4 = "1" then
      n16 <= n15;
    end if;
  end if;
end process;
n17 <= unsigned(signed(n6) * signed(n13));
n18 <= n17(34 downto 34) &
  n17(33 downto 33) &
  n17(32 downto 32) &
  n17(31 downto 31) &
  n17(30 downto 30) &
  n17(29 downto 29) &
  n17(28 downto 28) &
  n17(27 downto 27) &
  n17(26 downto 26) &
  n17(25 downto 25) &
  n17(24 downto 24) &
  n17(23 downto 23) &
  n17(22 downto 22) &
  n17(21 downto 21) &
  n17(20 downto 20) &
  n17(19 downto 19) &
  n17(18 downto 18) &
  n17(17 downto 17);
process (clock_c) begin
  if rising_edge(clock_c) then
    if i5 = "1" then
      n19 <= "000000000000000000";
    elsif i4 = "1" then
      n19 <= n18;
    end if;
  end if;
end process;
n20 <= n16 - n19;
process (clock_c) begin
  if rising_edge(clock_c) then
    if i5 = "1" then
      n21 <= "000000000000000000";
    elsif i4 = "1" then
      n21 <= n20;
    end if;
  end if;
end process;
n22 <= unsigned(signed(n5) * signed(n13));
n23 <= n22(34 downto 34) &
  n22(33 downto 33) &
  n22(32 downto 32) &
  n22(31 downto 31) &
  n22(30 downto 30) &
  n22(29 downto 29) &
  n22(28 downto 28) &
  n22(27 downto 27) &
  n22(26 downto 26) &
  n22(25 downto 25) &
  n22(24 downto 24) &
  n22(23 downto 23) &
  n22(22 downto 22) &
  n22(21 downto 21) &
  n22(20 downto 20) &
  n22(19 downto 19) &
  n22(18 downto 18) &
  n22(17 downto 17);
process (clock_c) begin
  if rising_edge(clock_c) then
    if i5 = "1" then
      n24 <= "000000000000000000";
    elsif i4 = "1" then
      n24 <= n23;
    end if;
  end if;
end process;
n25 <= unsigned(signed(n6) * signed(n12));
n26 <= n25(34 downto 34) &
  n25(33 downto 33) &
  n25(32 downto 32) &
  n25(31 downto 31) &
  n25(30 downto 30) &
  n25(29 downto 29) &
  n25(28 downto 28) &
  n25(27 downto 27) &
  n25(26 downto 26) &
  n25(25 downto 25) &
  n25(24 downto 24) &
  n25(23 downto 23) &
  n25(22 downto 22) &
  n25(21 downto 21) &
  n25(20 downto 20) &
  n25(19 downto 19) &
  n25(18 downto 18) &
  n25(17 downto 17);
process (clock_c) begin
  if rising_edge(clock_c) then
    if i5 = "1" then
      n27 <= "000000000000000000";
    elsif i4 = "1" then
      n27 <= n26;
    end if;
  end if;
end process;
n28 <= n24 + n27;
process (clock_c) begin
  if rising_edge(clock_c) then
    if i5 = "1" then
      n29 <= "000000000000000000";
    elsif i4 = "1" then
      n29 <= n28;
    end if;
  end if;
end process;
n30 <= n8 + n21;
n31 <= n10 + n29;
n32 <= n30 & n31;
process (clock_c) begin
  if rising_edge(clock_c) then
    if i5 = "1" then
      n33 <= "000000000000000000000000000000000000";
    elsif i4 = "1" then
      n33 <= n32;
    end if;
  end if;
end process;
n34 <= n8 - n21;
n35 <= n10 - n29;
n36 <= n34 & n35;
process (clock_c) begin
  if rising_edge(clock_c) then
    if i5 = "1" then
      n37 <= "000000000000000000000000000000000000";
    elsif i4 = "1" then
      n37 <= n36;
    end if;
  end if;
end process;
o2 <= n37;
o1 <= n33;
end architecture rtl;

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
entity cf_fft_256_18_18 is
port (
clock_c : in std_logic;
i1 : in  unsigned(71 downto 0);
i2 : in  unsigned(0 downto 0);
i3 : in  unsigned(5 downto 0);
i4 : in  unsigned(0 downto 0);
i5 : in  unsigned(0 downto 0);
i6 : in  unsigned(0 downto 0);
o1 : out unsigned(0 downto 0);
o2 : out unsigned(0 downto 0);
o3 : out unsigned(71 downto 0));
end entity cf_fft_256_18_18;
architecture rtl of cf_fft_256_18_18 is
signal n1 : unsigned(5 downto 0);
signal n2 : unsigned(5 downto 0);
signal n3 : unsigned(5 downto 0) := "000000";
signal n4 : unsigned(0 downto 0);
signal n5 : unsigned(0 downto 0) := "0";
signal n6 : unsigned(5 downto 0);
signal n7 : unsigned(0 downto 0);
signal n8 : unsigned(0 downto 0);
signal n9 : unsigned(71 downto 0);
signal n9a : unsigned(5 downto 0) := "000000";
type   n9mt is array (63 downto 0) of unsigned(71 downto 0);
signal n9m : n9mt;
signal n10 : unsigned(0 downto 0);
signal n11 : unsigned(71 downto 0);
signal n11a : unsigned(5 downto 0) := "000000";
type   n11mt is array (63 downto 0) of unsigned(71 downto 0);
signal n11m : n11mt;
signal n12 : unsigned(0 downto 0) := "0";
signal n13 : unsigned(71 downto 0);
signal n14 : unsigned(0 downto 0);
signal s15_1 : unsigned(0 downto 0);
component cf_fft_256_18_27 is
port (
clock_c : in std_logic;
i1 : in  unsigned(0 downto 0);
i2 : in  unsigned(0 downto 0);
i3 : in  unsigned(0 downto 0);
o1 : out unsigned(0 downto 0));
end component cf_fft_256_18_27;
begin
n1 <= "000001";
n2 <= n3 + n1;
process (clock_c) begin
  if rising_edge(clock_c) then
    if n14 = "1" then
      n3 <= "000000";
    elsif i5 = "1" then
      n3 <= n2;
    end if;
  end if;
end process;
n4 <= not s15_1;
process (clock_c) begin
  if rising_edge(clock_c) then
    if i6 = "1" then
      n5 <= "0";
    elsif i5 = "1" then
      n5 <= i2;
    end if;
  end if;
end process;
n6 <= "000000";
n7 <= "1" when n3 = n6 else "0";
n8 <= i4 and n4;
process (clock_c) begin
  if rising_edge(clock_c) then
    if i5 = "1" then
      if n8 = "1" then
        n9m(to_integer(i3)) <= i1;
      end if;
      n9a <= n3;
    end if;
  end if;
end process;
n9 <= n9m(to_integer(n9a));
n10 <= i4 and s15_1;
process (clock_c) begin
  if rising_edge(clock_c) then
    if i5 = "1" then
      if n10 = "1" then
        n11m(to_integer(i3)) <= i1;
      end if;
      n11a <= n3;
    end if;
  end if;
end process;
n11 <= n11m(to_integer(n11a));
process (clock_c) begin
  if rising_edge(clock_c) then
    if i6 = "1" then
      n12 <= "0";
    elsif i5 = "1" then
      n12 <= n4;
    end if;
  end if;
end process;
n13 <= n11 when n12 = "1" else n9;
n14 <= i2 or i6;
s15 : cf_fft_256_18_27 port map (clock_c, i2, i5, i6, s15_1);
o3 <= n13;
o2 <= n7;
o1 <= n5;
end architecture rtl;

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
entity cf_fft_256_18_17 is
port (
clock_c : in std_logic;
i1 : in  unsigned(71 downto 0);
i2 : in  unsigned(0 downto 0);
i3 : in  unsigned(5 downto 0);
i4 : in  unsigned(0 downto 0);
i5 : in  unsigned(0 downto 0);
i6 : in  unsigned(0 downto 0);
o1 : out unsigned(71 downto 0));
end entity cf_fft_256_18_17;
architecture rtl of cf_fft_256_18_17 is
signal n1 : unsigned(5 downto 0);
signal n2 : unsigned(5 downto 0);
signal n3 : unsigned(5 downto 0) := "000000";
signal n4 : unsigned(0 downto 0);
signal n5 : unsigned(0 downto 0);
signal n6 : unsigned(71 downto 0);
signal n6a : unsigned(5 downto 0) := "000000";
type   n6mt is array (63 downto 0) of unsigned(71 downto 0);
signal n6m : n6mt;
signal n7 : unsigned(0 downto 0);
signal n8 : unsigned(71 downto 0);
signal n8a : unsigned(5 downto 0) := "000000";
type   n8mt is array (63 downto 0) of unsigned(71 downto 0);
signal n8m : n8mt;
signal n9 : unsigned(0 downto 0) := "0";
signal n10 : unsigned(71 downto 0);
signal n11 : unsigned(0 downto 0);
signal s12_1 : unsigned(0 downto 0);
component cf_fft_256_18_27 is
port (
clock_c : in std_logic;
i1 : in  unsigned(0 downto 0);
i2 : in  unsigned(0 downto 0);
i3 : in  unsigned(0 downto 0);
o1 : out unsigned(0 downto 0));
end component cf_fft_256_18_27;
begin
n1 <= "000001";
n2 <= n3 + n1;
process (clock_c) begin
  if rising_edge(clock_c) then
    if n11 = "1" then
      n3 <= "000000";
    elsif i5 = "1" then
      n3 <= n2;
    end if;
  end if;
end process;
n4 <= not s12_1;
n5 <= i4 and n4;
process (clock_c) begin
  if rising_edge(clock_c) then
    if i5 = "1" then
      if n5 = "1" then
        n6m(to_integer(i3)) <= i1;
      end if;
      n6a <= n3;
    end if;
  end if;
end process;
n6 <= n6m(to_integer(n6a));
n7 <= i4 and s12_1;
process (clock_c) begin
  if rising_edge(clock_c) then
    if i5 = "1" then
      if n7 = "1" then
        n8m(to_integer(i3)) <= i1;
      end if;
      n8a <= n3;
    end if;
  end if;
end process;
n8 <= n8m(to_integer(n8a));
process (clock_c) begin
  if rising_edge(clock_c) then
    if i6 = "1" then
      n9 <= "0";
    elsif i5 = "1" then
      n9 <= n4;
    end if;
  end if;
end process;
n10 <= n8 when n9 = "1" else n6;
n11 <= i2 or i6;
s12 : cf_fft_256_18_27 port map (clock_c, i2, i5, i6, s12_1);
o1 <= n10;
end architecture rtl;

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
entity cf_fft_256_18_16 is
port (
clock_c : in std_logic;
i1 : in  unsigned(0 downto 0);
i2 : in  unsigned(35 downto 0);
i3 : in  unsigned(35 downto 0);
i4 : in  unsigned(0 downto 0);
i5 : in  unsigned(0 downto 0);
o1 : out unsigned(0 downto 0);
o2 : out unsigned(35 downto 0);
o3 : out unsigned(35 downto 0));
end entity cf_fft_256_18_16;
architecture rtl of cf_fft_256_18_16 is
signal n1 : unsigned(5 downto 0);
signal n2 : unsigned(71 downto 0);
signal n3 : unsigned(0 downto 0) := "0";
signal n4 : unsigned(0 downto 0) := "0";
signal n5 : unsigned(0 downto 0) := "0";
signal n6 : unsigned(0 downto 0) := "0";
signal n7 : unsigned(5 downto 0);
signal n8 : unsigned(5 downto 0) := "000000";
signal n9 : unsigned(5 downto 0) := "000000";
signal n10 : unsigned(5 downto 0) := "000000";
signal n11 : unsigned(5 downto 0) := "000000";
signal n12 : unsigned(0 downto 0);
signal n13 : unsigned(0 downto 0) := "0";
signal n14 : unsigned(0 downto 0) := "0";
signal n15 : unsigned(0 downto 0) := "0";
signal n16 : unsigned(0 downto 0) := "0";
signal n17 : unsigned(0 downto 0);
signal n18 : unsigned(1 downto 0);
signal n19 : unsigned(35 downto 0);
signal n20 : unsigned(35 downto 0);
signal n21 : unsigned(35 downto 0);
signal n22 : unsigned(35 downto 0);
signal n23 : unsigned(35 downto 0);
signal n24 : unsigned(35 downto 0);
signal s25_1 : unsigned(0 downto 0);
signal s26_1 : unsigned(35 downto 0);
signal s26_2 : unsigned(35 downto 0);
signal s27_1 : unsigned(6 downto 0);
signal s27_2 : unsigned(0 downto 0);
signal s28_1 : unsigned(0 downto 0);
signal s28_2 : unsigned(0 downto 0);
signal s28_3 : unsigned(71 downto 0);
signal s29_1 : unsigned(71 downto 0);
component cf_fft_256_18_30 is
port (
clock_c : in std_logic;
i1 : in  unsigned(1 downto 0);
i2 : in  unsigned(0 downto 0);
i3 : in  unsigned(0 downto 0);
o1 : out unsigned(0 downto 0));
end component cf_fft_256_18_30;
component cf_fft_256_18_19 is
port (
clock_c : in std_logic;
i1 : in  unsigned(35 downto 0);
i2 : in  unsigned(35 downto 0);
i3 : in  unsigned(5 downto 0);
i4 : in  unsigned(0 downto 0);
i5 : in  unsigned(0 downto 0);
o1 : out unsigned(35 downto 0);
o2 : out unsigned(35 downto 0));
end component cf_fft_256_18_19;
component cf_fft_256_18_21 is
port (
clock_c : in std_logic;
i1 : in  unsigned(0 downto 0);
i2 : in  unsigned(0 downto 0);
i3 : in  unsigned(0 downto 0);
o1 : out unsigned(6 downto 0);
o2 : out unsigned(0 downto 0));
end component cf_fft_256_18_21;
component cf_fft_256_18_18 is
port (
clock_c : in std_logic;
i1 : in  unsigned(71 downto 0);
i2 : in  unsigned(0 downto 0);
i3 : in  unsigned(5 downto 0);
i4 : in  unsigned(0 downto 0);
i5 : in  unsigned(0 downto 0);
i6 : in  unsigned(0 downto 0);
o1 : out unsigned(0 downto 0);
o2 : out unsigned(0 downto 0);
o3 : out unsigned(71 downto 0));
end component cf_fft_256_18_18;
component cf_fft_256_18_17 is
port (
clock_c : in std_logic;
i1 : in  unsigned(71 downto 0);
i2 : in  unsigned(0 downto 0);
i3 : in  unsigned(5 downto 0);
i4 : in  unsigned(0 downto 0);
i5 : in  unsigned(0 downto 0);
i6 : in  unsigned(0 downto 0);
o1 : out unsigned(71 downto 0));
end component cf_fft_256_18_17;
begin
n1 <= s27_1(6 downto 6) &
  s27_1(5 downto 5) &
  s27_1(4 downto 4) &
  s27_1(3 downto 3) &
  s27_1(2 downto 2) &
  s27_1(1 downto 1);
n2 <= s26_1 & s26_2;
process (clock_c) begin
  if rising_edge(clock_c) then
    if i5 = "1" then
      n3 <= "0";
    elsif i4 = "1" then
      n3 <= s27_2;
    end if;
  end if;
end process;
process (clock_c) begin
  if rising_edge(clock_c) then
    if i5 = "1" then
      n4 <= "0";
    elsif i4 = "1" then
      n4 <= n3;
    end if;
  end if;
end process;
process (clock_c) begin
  if rising_edge(clock_c) then
    if i5 = "1" then
      n5 <= "0";
    elsif i4 = "1" then
      n5 <= n4;
    end if;
  end if;
end process;
process (clock_c) begin
  if rising_edge(clock_c) then
    if i5 = "1" then
      n6 <= "0";
    elsif i4 = "1" then
      n6 <= n5;
    end if;
  end if;
end process;
n7 <= s27_1(6 downto 6) &
  s27_1(5 downto 5) &
  s27_1(4 downto 4) &
  s27_1(3 downto 3) &
  s27_1(2 downto 2) &
  s27_1(1 downto 1);
process (clock_c) begin
  if rising_edge(clock_c) then
    if i5 = "1" then
      n8 <= "000000";
    elsif i4 = "1" then
      n8 <= n7;
    end if;
  end if;
end process;
process (clock_c) begin
  if rising_edge(clock_c) then
    if i5 = "1" then
      n9 <= "000000";
    elsif i4 = "1" then
      n9 <= n8;
    end if;
  end if;
end process;
process (clock_c) begin
  if rising_edge(clock_c) then
    if i5 = "1" then
      n10 <= "000000";
    elsif i4 = "1" then
      n10 <= n9;
    end if;
  end if;
end process;
process (clock_c) begin
  if rising_edge(clock_c) then
    if i5 = "1" then
      n11 <= "000000";
    elsif i4 = "1" then
      n11 <= n10;
    end if;
  end if;
end process;
n12 <= s27_1(0 downto 0);
process (clock_c) begin
  if rising_edge(clock_c) then
    if i5 = "1" then
      n13 <= "0";
    elsif i4 = "1" then
      n13 <= n12;
    end if;
  end if;
end process;
process (clock_c) begin
  if rising_edge(clock_c) then
    if i5 = "1" then
      n14 <= "0";
    elsif i4 = "1" then
      n14 <= n13;
    end if;
  end if;
end process;
process (clock_c) begin
  if rising_edge(clock_c) then
    if i5 = "1" then
      n15 <= "0";
    elsif i4 = "1" then
      n15 <= n14;
    end if;
  end if;
end process;
process (clock_c) begin
  if rising_edge(clock_c) then
    if i5 = "1" then
      n16 <= "0";
    elsif i4 = "1" then
      n16 <= n15;
    end if;
  end if;
end process;
n17 <= not n16;
n18 <= s28_2 & s28_1;
n19 <= s28_3(71 downto 71) &
  s28_3(70 downto 70) &
  s28_3(69 downto 69) &
  s28_3(68 downto 68) &
  s28_3(67 downto 67) &
  s28_3(66 downto 66) &
  s28_3(65 downto 65) &
  s28_3(64 downto 64) &
  s28_3(63 downto 63) &
  s28_3(62 downto 62) &
  s28_3(61 downto 61) &
  s28_3(60 downto 60) &
  s28_3(59 downto 59) &
  s28_3(58 downto 58) &
  s28_3(57 downto 57) &
  s28_3(56 downto 56) &
  s28_3(55 downto 55) &
  s28_3(54 downto 54) &
  s28_3(53 downto 53) &
  s28_3(52 downto 52) &
  s28_3(51 downto 51) &
  s28_3(50 downto 50) &
  s28_3(49 downto 49) &
  s28_3(48 downto 48) &
  s28_3(47 downto 47) &
  s28_3(46 downto 46) &
  s28_3(45 downto 45) &
  s28_3(44 downto 44) &
  s28_3(43 downto 43) &
  s28_3(42 downto 42) &
  s28_3(41 downto 41) &
  s28_3(40 downto 40) &
  s28_3(39 downto 39) &
  s28_3(38 downto 38) &
  s28_3(37 downto 37) &
  s28_3(36 downto 36);
n20 <= s28_3(35 downto 35) &
  s28_3(34 downto 34) &
  s28_3(33 downto 33) &
  s28_3(32 downto 32) &
  s28_3(31 downto 31) &
  s28_3(30 downto 30) &
  s28_3(29 downto 29) &
  s28_3(28 downto 28) &
  s28_3(27 downto 27) &
  s28_3(26 downto 26) &
  s28_3(25 downto 25) &
  s28_3(24 downto 24) &
  s28_3(23 downto 23) &
  s28_3(22 downto 22) &
  s28_3(21 downto 21) &
  s28_3(20 downto 20) &
  s28_3(19 downto 19) &
  s28_3(18 downto 18) &
  s28_3(17 downto 17) &
  s28_3(16 downto 16) &
  s28_3(15 downto 15) &
  s28_3(14 downto 14) &
  s28_3(13 downto 13) &
  s28_3(12 downto 12) &
  s28_3(11 downto 11) &
  s28_3(10 downto 10) &
  s28_3(9 downto 9) &
  s28_3(8 downto 8) &
  s28_3(7 downto 7) &
  s28_3(6 downto 6) &
  s28_3(5 downto 5) &
  s28_3(4 downto 4) &
  s28_3(3 downto 3) &
  s28_3(2 downto 2) &
  s28_3(1 downto 1) &
  s28_3(0 downto 0);
n21 <= s29_1(71 downto 71) &
  s29_1(70 downto 70) &
  s29_1(69 downto 69) &
  s29_1(68 downto 68) &
  s29_1(67 downto 67) &
  s29_1(66 downto 66) &
  s29_1(65 downto 65) &
  s29_1(64 downto 64) &
  s29_1(63 downto 63) &
  s29_1(62 downto 62) &
  s29_1(61 downto 61) &
  s29_1(60 downto 60) &
  s29_1(59 downto 59) &
  s29_1(58 downto 58) &
  s29_1(57 downto 57) &
  s29_1(56 downto 56) &
  s29_1(55 downto 55) &
  s29_1(54 downto 54) &
  s29_1(53 downto 53) &
  s29_1(52 downto 52) &
  s29_1(51 downto 51) &
  s29_1(50 downto 50) &
  s29_1(49 downto 49) &
  s29_1(48 downto 48) &
  s29_1(47 downto 47) &
  s29_1(46 downto 46) &
  s29_1(45 downto 45) &
  s29_1(44 downto 44) &
  s29_1(43 downto 43) &
  s29_1(42 downto 42) &
  s29_1(41 downto 41) &
  s29_1(40 downto 40) &
  s29_1(39 downto 39) &
  s29_1(38 downto 38) &
  s29_1(37 downto 37) &
  s29_1(36 downto 36);
n22 <= s29_1(35 downto 35) &
  s29_1(34 downto 34) &
  s29_1(33 downto 33) &
  s29_1(32 downto 32) &
  s29_1(31 downto 31) &
  s29_1(30 downto 30) &
  s29_1(29 downto 29) &
  s29_1(28 downto 28) &
  s29_1(27 downto 27) &
  s29_1(26 downto 26) &
  s29_1(25 downto 25) &
  s29_1(24 downto 24) &
  s29_1(23 downto 23) &
  s29_1(22 downto 22) &
  s29_1(21 downto 21) &
  s29_1(20 downto 20) &
  s29_1(19 downto 19) &
  s29_1(18 downto 18) &
  s29_1(17 downto 17) &
  s29_1(16 downto 16) &
  s29_1(15 downto 15) &
  s29_1(14 downto 14) &
  s29_1(13 downto 13) &
  s29_1(12 downto 12) &
  s29_1(11 downto 11) &
  s29_1(10 downto 10) &
  s29_1(9 downto 9) &
  s29_1(8 downto 8) &
  s29_1(7 downto 7) &
  s29_1(6 downto 6) &
  s29_1(5 downto 5) &
  s29_1(4 downto 4) &
  s29_1(3 downto 3) &
  s29_1(2 downto 2) &
  s29_1(1 downto 1) &
  s29_1(0 downto 0);
n23 <= n20 when s25_1 = "1" else n19;
n24 <= n22 when s25_1 = "1" else n21;
s25 : cf_fft_256_18_30 port map (clock_c, n18, i4, i5, s25_1);
s26 : cf_fft_256_18_19 port map (clock_c, i2, i3, n1, i4, i5, s26_1, s26_2);
s27 : cf_fft_256_18_21 port map (clock_c, i1, i4, i5, s27_1, s27_2);
s28 : cf_fft_256_18_18 port map (clock_c, n2, n6, n11, n17, i4, i5, s28_1, s28_2, s28_3);
s29 : cf_fft_256_18_17 port map (clock_c, n2, n6, n11, n16, i4, i5, s29_1);
o3 <= n24;
o2 <= n23;
o1 <= s28_1;
end architecture rtl;

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
entity cf_fft_256_18_15 is
port (
clock_c : in std_logic;
i1 : in  unsigned(35 downto 0);
i2 : in  unsigned(35 downto 0);
i3 : in  unsigned(6 downto 0);
i4 : in  unsigned(0 downto 0);
i5 : in  unsigned(0 downto 0);
o1 : out unsigned(35 downto 0);
o2 : out unsigned(35 downto 0));
end entity cf_fft_256_18_15;
architecture rtl of cf_fft_256_18_15 is
signal n1 : unsigned(35 downto 0) := "000000000000000000000000000000000000";
signal n2 : unsigned(17 downto 0);
signal n3 : unsigned(17 downto 0);
signal n4 : unsigned(35 downto 0) := "000000000000000000000000000000000000";
signal n5 : unsigned(17 downto 0);
signal n6 : unsigned(17 downto 0);
signal n7 : unsigned(17 downto 0) := "000000000000000000";
signal n8 : unsigned(17 downto 0) := "000000000000000000";
signal n9 : unsigned(17 downto 0) := "000000000000000000";
signal n10 : unsigned(17 downto 0) := "000000000000000000";
signal n11 : unsigned(35 downto 0) := "000000000000000000000000000000000000";
signal n12 : unsigned(17 downto 0);
signal n13 : unsigned(17 downto 0);
signal n14 : unsigned(35 downto 0);
signal n15 : unsigned(17 downto 0);
signal n16 : unsigned(17 downto 0) := "000000000000000000";
signal n17 : unsigned(35 downto 0);
signal n18 : unsigned(17 downto 0);
signal n19 : unsigned(17 downto 0) := "000000000000000000";
signal n20 : unsigned(17 downto 0);
signal n21 : unsigned(17 downto 0) := "000000000000000000";
signal n22 : unsigned(35 downto 0);
signal n23 : unsigned(17 downto 0);
signal n24 : unsigned(17 downto 0) := "000000000000000000";
signal n25 : unsigned(35 downto 0);
signal n26 : unsigned(17 downto 0);
signal n27 : unsigned(17 downto 0) := "000000000000000000";
signal n28 : unsigned(17 downto 0);
signal n29 : unsigned(17 downto 0) := "000000000000000000";
signal n30 : unsigned(17 downto 0);
signal n31 : unsigned(17 downto 0);
signal n32 : unsigned(35 downto 0);
signal n33 : unsigned(35 downto 0) := "000000000000000000000000000000000000";
signal n34 : unsigned(17 downto 0);
signal n35 : unsigned(17 downto 0);
signal n36 : unsigned(35 downto 0);
signal n37 : unsigned(35 downto 0) := "000000000000000000000000000000000000";
begin
process (clock_c) begin
  if rising_edge(clock_c) then
    if i5 = "1" then
      n1 <= "000000000000000000000000000000000000";
    elsif i4 = "1" then
      n1 <= i1;
    end if;
  end if;
end process;
n2 <= n1(35 downto 35) &
  n1(34 downto 34) &
  n1(33 downto 33) &
  n1(32 downto 32) &
  n1(31 downto 31) &
  n1(30 downto 30) &
  n1(29 downto 29) &
  n1(28 downto 28) &
  n1(27 downto 27) &
  n1(26 downto 26) &
  n1(25 downto 25) &
  n1(24 downto 24) &
  n1(23 downto 23) &
  n1(22 downto 22) &
  n1(21 downto 21) &
  n1(20 downto 20) &
  n1(19 downto 19) &
  n1(18 downto 18);
n3 <= n1(17 downto 17) &
  n1(16 downto 16) &
  n1(15 downto 15) &
  n1(14 downto 14) &
  n1(13 downto 13) &
  n1(12 downto 12) &
  n1(11 downto 11) &
  n1(10 downto 10) &
  n1(9 downto 9) &
  n1(8 downto 8) &
  n1(7 downto 7) &
  n1(6 downto 6) &
  n1(5 downto 5) &
  n1(4 downto 4) &
  n1(3 downto 3) &
  n1(2 downto 2) &
  n1(1 downto 1) &
  n1(0 downto 0);
process (clock_c) begin
  if rising_edge(clock_c) then
    if i5 = "1" then
      n4 <= "000000000000000000000000000000000000";
    elsif i4 = "1" then
      n4 <= i2;
    end if;
  end if;
end process;
n5 <= n4(35 downto 35) &
  n4(34 downto 34) &
  n4(33 downto 33) &
  n4(32 downto 32) &
  n4(31 downto 31) &
  n4(30 downto 30) &
  n4(29 downto 29) &
  n4(28 downto 28) &
  n4(27 downto 27) &
  n4(26 downto 26) &
  n4(25 downto 25) &
  n4(24 downto 24) &
  n4(23 downto 23) &
  n4(22 downto 22) &
  n4(21 downto 21) &
  n4(20 downto 20) &
  n4(19 downto 19) &
  n4(18 downto 18);
n6 <= n4(17 downto 17) &
  n4(16 downto 16) &
  n4(15 downto 15) &
  n4(14 downto 14) &
  n4(13 downto 13) &
  n4(12 downto 12) &
  n4(11 downto 11) &
  n4(10 downto 10) &
  n4(9 downto 9) &
  n4(8 downto 8) &
  n4(7 downto 7) &
  n4(6 downto 6) &
  n4(5 downto 5) &
  n4(4 downto 4) &
  n4(3 downto 3) &
  n4(2 downto 2) &
  n4(1 downto 1) &
  n4(0 downto 0);
process (clock_c) begin
  if rising_edge(clock_c) then
    if i5 = "1" then
      n7 <= "000000000000000000";
    elsif i4 = "1" then
      n7 <= n2;
    end if;
  end if;
end process;
process (clock_c) begin
  if rising_edge(clock_c) then
    if i5 = "1" then
      n8 <= "000000000000000000";
    elsif i4 = "1" then
      n8 <= n7;
    end if;
  end if;
end process;
process (clock_c) begin
  if rising_edge(clock_c) then
    if i5 = "1" then
      n9 <= "000000000000000000";
    elsif i4 = "1" then
      n9 <= n3;
    end if;
  end if;
end process;
process (clock_c) begin
  if rising_edge(clock_c) then
    if i5 = "1" then
      n10 <= "000000000000000000";
    elsif i4 = "1" then
      n10 <= n9;
    end if;
  end if;
end process;
process (clock_c) begin
  if rising_edge(clock_c) then 
    if i4 = "1" then
      case i3 is
        when "0000000" => n11 <= "011111111111111111000000000000000000";
        when "0000001" => n11 <= "011111111111011000111111001101101111";
        when "0000010" => n11 <= "011111111101100010111110011011100000";
        when "0000011" => n11 <= "011111111010011100111101101001010101";
        when "0000100" => n11 <= "011111110110001000111100110111010000";
        when "0000101" => n11 <= "011111110000100110111100000101010011";
        when "0000110" => n11 <= "011111101001110101111011010011011111";
        when "0000111" => n11 <= "011111100001110110111010100001110111";
        when "0001000" => n11 <= "011111011000101001111001110000011101";
        when "0001001" => n11 <= "011111001110001111111000111111010001";
        when "0001010" => n11 <= "011111000010100111111000001110011000";
        when "0001011" => n11 <= "011110110101110100110111011101110001";
        when "0001100" => n11 <= "011110100111110100110110101101011111";
        when "0001101" => n11 <= "011110011000101000110101111101100101";
        when "0001110" => n11 <= "011110001000010010110101001110000011";
        when "0001111" => n11 <= "011101110110110001110100011110111011";
        when "0010000" => n11 <= "011101100100000110110011110000010000";
        when "0010001" => n11 <= "011101010000010011110011000010000100";
        when "0010010" => n11 <= "011100111011010111110010010100010111";
        when "0010011" => n11 <= "011100100101010100110001100111001100";
        when "0010100" => n11 <= "011100001110001011110000111010100101";
        when "0010101" => n11 <= "011011110101111100110000001110100010";
        when "0010110" => n11 <= "011011011100101000101111100011000111";
        when "0010111" => n11 <= "011011000010010000101110111000010100";
        when "0011000" => n11 <= "011010100110110110101110001110001100";
        when "0011001" => n11 <= "011010001010011010101101100100101111";
        when "0011010" => n11 <= "011001101100111110101100111100000000";
        when "0011011" => n11 <= "011001001110100010101100010100000000";
        when "0011100" => n11 <= "011000101111001000101011101100110000";
        when "0011101" => n11 <= "011000001110110000101011000110010011";
        when "0011110" => n11 <= "010111101101011101101010100000101001";
        when "0011111" => n11 <= "010111001011010000101001111011110100";
        when "0100000" => n11 <= "010110101000001001101001010111110110";
        when "0100001" => n11 <= "010110000100001011101000110100101111";
        when "0100010" => n11 <= "010101011111010110101000010010100010";
        when "0100011" => n11 <= "010100111001101100100111110001001111";
        when "0100100" => n11 <= "010100010011001111100111010000110111";
        when "0100101" => n11 <= "010011101011111111100110110001011101";
        when "0100110" => n11 <= "010011000011111111100110010011000001";
        when "0100111" => n11 <= "010010011011010000100101110101100101";
        when "0101000" => n11 <= "010001110001110011100101011001001001";
        when "0101001" => n11 <= "010001000111101011100100111101101111";
        when "0101010" => n11 <= "010000011100111000100100100011010111";
        when "0101011" => n11 <= "001111110001011101100100001010000011";
        when "0101100" => n11 <= "001111000101011010100011110001110100";
        when "0101101" => n11 <= "001110011000110011100011011010101011";
        when "0101110" => n11 <= "001101101011101000100011000100101000";
        when "0101111" => n11 <= "001100111101111011100010101111101100";
        when "0110000" => n11 <= "001100001111101111100010011011111001";
        when "0110001" => n11 <= "001011100001000100100010001001001110";
        when "0110010" => n11 <= "001010110001111100100001110111101101";
        when "0110011" => n11 <= "001010000010011010100001100111010111";
        when "0110100" => n11 <= "001001010010100000100001011000001011";
        when "0110101" => n11 <= "001000100010001110100001001010001011";
        when "0110110" => n11 <= "000111110001100111100000111101011000";
        when "0110111" => n11 <= "000111000000101110100000110001110000";
        when "0111000" => n11 <= "000110001111100010100000100111010110";
        when "0111001" => n11 <= "000101011110001000100000011110001001";
        when "0111010" => n11 <= "000100101100100000100000010110001010";
        when "0111011" => n11 <= "000011111010101100100000001111011001";
        when "0111100" => n11 <= "000011001000101111100000001001110111";
        when "0111101" => n11 <= "000010010110101010100000000101100011";
        when "0111110" => n11 <= "000001100100011111100000000010011101";
        when "0111111" => n11 <= "000000110010010000100000000000100111";
        when "1000000" => n11 <= "000000000000000000100000000000000000";
        when "1000001" => n11 <= "111111001101101111100000000000100111";
        when "1000010" => n11 <= "111110011011100000100000000010011101";
        when "1000011" => n11 <= "111101101001010101100000000101100011";
        when "1000100" => n11 <= "111100110111010000100000001001110111";
        when "1000101" => n11 <= "111100000101010011100000001111011001";
        when "1000110" => n11 <= "111011010011011111100000010110001010";
        when "1000111" => n11 <= "111010100001110111100000011110001001";
        when "1001000" => n11 <= "111001110000011101100000100111010110";
        when "1001001" => n11 <= "111000111111010001100000110001110000";
        when "1001010" => n11 <= "111000001110011000100000111101011000";
        when "1001011" => n11 <= "110111011101110001100001001010001011";
        when "1001100" => n11 <= "110110101101011111100001011000001011";
        when "1001101" => n11 <= "110101111101100101100001100111010111";
        when "1001110" => n11 <= "110101001110000011100001110111101101";
        when "1001111" => n11 <= "110100011110111011100010001001001110";
        when "1010000" => n11 <= "110011110000010000100010011011111001";
        when "1010001" => n11 <= "110011000010000100100010101111101100";
        when "1010010" => n11 <= "110010010100010111100011000100101000";
        when "1010011" => n11 <= "110001100111001100100011011010101011";
        when "1010100" => n11 <= "110000111010100101100011110001110100";
        when "1010101" => n11 <= "110000001110100010100100001010000011";
        when "1010110" => n11 <= "101111100011000111100100100011010111";
        when "1010111" => n11 <= "101110111000010100100100111101101111";
        when "1011000" => n11 <= "101110001110001100100101011001001001";
        when "1011001" => n11 <= "101101100100101111100101110101100101";
        when "1011010" => n11 <= "101100111100000000100110010011000001";
        when "1011011" => n11 <= "101100010100000000100110110001011101";
        when "1011100" => n11 <= "101011101100110000100111010000110111";
        when "1011101" => n11 <= "101011000110010011100111110001001111";
        when "1011110" => n11 <= "101010100000101001101000010010100010";
        when "1011111" => n11 <= "101001111011110100101000110100101111";
        when "1100000" => n11 <= "101001010111110110101001010111110110";
        when "1100001" => n11 <= "101000110100101111101001111011110100";
        when "1100010" => n11 <= "101000010010100010101010100000101001";
        when "1100011" => n11 <= "100111110001001111101011000110010011";
        when "1100100" => n11 <= "100111010000110111101011101100110000";
        when "1100101" => n11 <= "100110110001011101101100010100000000";
        when "1100110" => n11 <= "100110010011000001101100111100000000";
        when "1100111" => n11 <= "100101110101100101101101100100101111";
        when "1101000" => n11 <= "100101011001001001101110001110001100";
        when "1101001" => n11 <= "100100111101101111101110111000010100";
        when "1101010" => n11 <= "100100100011010111101111100011000111";
        when "1101011" => n11 <= "100100001010000011110000001110100010";
        when "1101100" => n11 <= "100011110001110100110000111010100101";
        when "1101101" => n11 <= "100011011010101011110001100111001100";
        when "1101110" => n11 <= "100011000100101000110010010100010111";
        when "1101111" => n11 <= "100010101111101100110011000010000100";
        when "1110000" => n11 <= "100010011011111001110011110000010000";
        when "1110001" => n11 <= "100010001001001110110100011110111011";
        when "1110010" => n11 <= "100001110111101101110101001110000011";
        when "1110011" => n11 <= "100001100111010111110101111101100101";
        when "1110100" => n11 <= "100001011000001011110110101101011111";
        when "1110101" => n11 <= "100001001010001011110111011101110001";
        when "1110110" => n11 <= "100000111101011000111000001110011000";
        when "1110111" => n11 <= "100000110001110000111000111111010001";
        when "1111000" => n11 <= "100000100111010110111001110000011101";
        when "1111001" => n11 <= "100000011110001001111010100001110111";
        when "1111010" => n11 <= "100000010110001010111011010011011111";
        when "1111011" => n11 <= "100000001111011001111100000101010011";
        when "1111100" => n11 <= "100000001001110111111100110111010000";
        when "1111101" => n11 <= "100000000101100011111101101001010101";
        when "1111110" => n11 <= "100000000010011101111110011011100000";
        when "1111111" => n11 <= "100000000000100111111111001101101111";
        when others => n11 <= "XXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX";
      end case;
    end if;
  end if;
end process;
n12 <= n11(35 downto 35) &
  n11(34 downto 34) &
  n11(33 downto 33) &
  n11(32 downto 32) &
  n11(31 downto 31) &
  n11(30 downto 30) &
  n11(29 downto 29) &
  n11(28 downto 28) &
  n11(27 downto 27) &
  n11(26 downto 26) &
  n11(25 downto 25) &
  n11(24 downto 24) &
  n11(23 downto 23) &
  n11(22 downto 22) &
  n11(21 downto 21) &
  n11(20 downto 20) &
  n11(19 downto 19) &
  n11(18 downto 18);
n13 <= n11(17 downto 17) &
  n11(16 downto 16) &
  n11(15 downto 15) &
  n11(14 downto 14) &
  n11(13 downto 13) &
  n11(12 downto 12) &
  n11(11 downto 11) &
  n11(10 downto 10) &
  n11(9 downto 9) &
  n11(8 downto 8) &
  n11(7 downto 7) &
  n11(6 downto 6) &
  n11(5 downto 5) &
  n11(4 downto 4) &
  n11(3 downto 3) &
  n11(2 downto 2) &
  n11(1 downto 1) &
  n11(0 downto 0);
n14 <= unsigned(signed(n5) * signed(n12));
n15 <= n14(34 downto 34) &
  n14(33 downto 33) &
  n14(32 downto 32) &
  n14(31 downto 31) &
  n14(30 downto 30) &
  n14(29 downto 29) &
  n14(28 downto 28) &
  n14(27 downto 27) &
  n14(26 downto 26) &
  n14(25 downto 25) &
  n14(24 downto 24) &
  n14(23 downto 23) &
  n14(22 downto 22) &
  n14(21 downto 21) &
  n14(20 downto 20) &
  n14(19 downto 19) &
  n14(18 downto 18) &
  n14(17 downto 17);
process (clock_c) begin
  if rising_edge(clock_c) then
    if i5 = "1" then
      n16 <= "000000000000000000";
    elsif i4 = "1" then
      n16 <= n15;
    end if;
  end if;
end process;
n17 <= unsigned(signed(n6) * signed(n13));
n18 <= n17(34 downto 34) &
  n17(33 downto 33) &
  n17(32 downto 32) &
  n17(31 downto 31) &
  n17(30 downto 30) &
  n17(29 downto 29) &
  n17(28 downto 28) &
  n17(27 downto 27) &
  n17(26 downto 26) &
  n17(25 downto 25) &
  n17(24 downto 24) &
  n17(23 downto 23) &
  n17(22 downto 22) &
  n17(21 downto 21) &
  n17(20 downto 20) &
  n17(19 downto 19) &
  n17(18 downto 18) &
  n17(17 downto 17);
process (clock_c) begin
  if rising_edge(clock_c) then
    if i5 = "1" then
      n19 <= "000000000000000000";
    elsif i4 = "1" then
      n19 <= n18;
    end if;
  end if;
end process;
n20 <= n16 - n19;
process (clock_c) begin
  if rising_edge(clock_c) then
    if i5 = "1" then
      n21 <= "000000000000000000";
    elsif i4 = "1" then
      n21 <= n20;
    end if;
  end if;
end process;
n22 <= unsigned(signed(n5) * signed(n13));
n23 <= n22(34 downto 34) &
  n22(33 downto 33) &
  n22(32 downto 32) &
  n22(31 downto 31) &
  n22(30 downto 30) &
  n22(29 downto 29) &
  n22(28 downto 28) &
  n22(27 downto 27) &
  n22(26 downto 26) &
  n22(25 downto 25) &
  n22(24 downto 24) &
  n22(23 downto 23) &
  n22(22 downto 22) &
  n22(21 downto 21) &
  n22(20 downto 20) &
  n22(19 downto 19) &
  n22(18 downto 18) &
  n22(17 downto 17);
process (clock_c) begin
  if rising_edge(clock_c) then
    if i5 = "1" then
      n24 <= "000000000000000000";
    elsif i4 = "1" then
      n24 <= n23;
    end if;
  end if;
end process;
n25 <= unsigned(signed(n6) * signed(n12));
n26 <= n25(34 downto 34) &
  n25(33 downto 33) &
  n25(32 downto 32) &
  n25(31 downto 31) &
  n25(30 downto 30) &
  n25(29 downto 29) &
  n25(28 downto 28) &
  n25(27 downto 27) &
  n25(26 downto 26) &
  n25(25 downto 25) &
  n25(24 downto 24) &
  n25(23 downto 23) &
  n25(22 downto 22) &
  n25(21 downto 21) &
  n25(20 downto 20) &
  n25(19 downto 19) &
  n25(18 downto 18) &
  n25(17 downto 17);
process (clock_c) begin
  if rising_edge(clock_c) then
    if i5 = "1" then
      n27 <= "000000000000000000";
    elsif i4 = "1" then
      n27 <= n26;
    end if;
  end if;
end process;
n28 <= n24 + n27;
process (clock_c) begin
  if rising_edge(clock_c) then
    if i5 = "1" then
      n29 <= "000000000000000000";
    elsif i4 = "1" then
      n29 <= n28;
    end if;
  end if;
end process;
n30 <= n8 + n21;
n31 <= n10 + n29;
n32 <= n30 & n31;
process (clock_c) begin
  if rising_edge(clock_c) then
    if i5 = "1" then
      n33 <= "000000000000000000000000000000000000";
    elsif i4 = "1" then
      n33 <= n32;
    end if;
  end if;
end process;
n34 <= n8 - n21;
n35 <= n10 - n29;
n36 <= n34 & n35;
process (clock_c) begin
  if rising_edge(clock_c) then
    if i5 = "1" then
      n37 <= "000000000000000000000000000000000000";
    elsif i4 = "1" then
      n37 <= n36;
    end if;
  end if;
end process;
o2 <= n37;
o1 <= n33;
end architecture rtl;

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
entity cf_fft_256_18_14 is
port (
clock_c : in std_logic;
i1 : in  unsigned(0 downto 0);
i2 : in  unsigned(35 downto 0);
i3 : in  unsigned(35 downto 0);
i4 : in  unsigned(0 downto 0);
i5 : in  unsigned(0 downto 0);
o1 : out unsigned(0 downto 0);
o2 : out unsigned(35 downto 0);
o3 : out unsigned(35 downto 0));
end entity cf_fft_256_18_14;
architecture rtl of cf_fft_256_18_14 is
signal n1 : unsigned(6 downto 0);
signal n2 : unsigned(71 downto 0);
signal n3 : unsigned(0 downto 0) := "0";
signal n4 : unsigned(0 downto 0) := "0";
signal n5 : unsigned(0 downto 0) := "0";
signal n6 : unsigned(0 downto 0) := "0";
signal n7 : unsigned(5 downto 0);
signal n8 : unsigned(5 downto 0) := "000000";
signal n9 : unsigned(5 downto 0) := "000000";
signal n10 : unsigned(5 downto 0) := "000000";
signal n11 : unsigned(5 downto 0) := "000000";
signal n12 : unsigned(0 downto 0);
signal n13 : unsigned(0 downto 0) := "0";
signal n14 : unsigned(0 downto 0) := "0";
signal n15 : unsigned(0 downto 0) := "0";
signal n16 : unsigned(0 downto 0) := "0";
signal n17 : unsigned(0 downto 0);
signal n18 : unsigned(1 downto 0);
signal n19 : unsigned(35 downto 0);
signal n20 : unsigned(35 downto 0);
signal n21 : unsigned(35 downto 0);
signal n22 : unsigned(35 downto 0);
signal n23 : unsigned(35 downto 0);
signal n24 : unsigned(35 downto 0);
signal s25_1 : unsigned(35 downto 0);
signal s25_2 : unsigned(35 downto 0);
signal s26_1 : unsigned(0 downto 0);
signal s27_1 : unsigned(6 downto 0);
signal s27_2 : unsigned(0 downto 0);
signal s28_1 : unsigned(71 downto 0);
signal s29_1 : unsigned(0 downto 0);
signal s29_2 : unsigned(0 downto 0);
signal s29_3 : unsigned(71 downto 0);
component cf_fft_256_18_15 is
port (
clock_c : in std_logic;
i1 : in  unsigned(35 downto 0);
i2 : in  unsigned(35 downto 0);
i3 : in  unsigned(6 downto 0);
i4 : in  unsigned(0 downto 0);
i5 : in  unsigned(0 downto 0);
o1 : out unsigned(35 downto 0);
o2 : out unsigned(35 downto 0));
end component cf_fft_256_18_15;
component cf_fft_256_18_30 is
port (
clock_c : in std_logic;
i1 : in  unsigned(1 downto 0);
i2 : in  unsigned(0 downto 0);
i3 : in  unsigned(0 downto 0);
o1 : out unsigned(0 downto 0));
end component cf_fft_256_18_30;
component cf_fft_256_18_21 is
port (
clock_c : in std_logic;
i1 : in  unsigned(0 downto 0);
i2 : in  unsigned(0 downto 0);
i3 : in  unsigned(0 downto 0);
o1 : out unsigned(6 downto 0);
o2 : out unsigned(0 downto 0));
end component cf_fft_256_18_21;
component cf_fft_256_18_17 is
port (
clock_c : in std_logic;
i1 : in  unsigned(71 downto 0);
i2 : in  unsigned(0 downto 0);
i3 : in  unsigned(5 downto 0);
i4 : in  unsigned(0 downto 0);
i5 : in  unsigned(0 downto 0);
i6 : in  unsigned(0 downto 0);
o1 : out unsigned(71 downto 0));
end component cf_fft_256_18_17;
component cf_fft_256_18_18 is
port (
clock_c : in std_logic;
i1 : in  unsigned(71 downto 0);
i2 : in  unsigned(0 downto 0);
i3 : in  unsigned(5 downto 0);
i4 : in  unsigned(0 downto 0);
i5 : in  unsigned(0 downto 0);
i6 : in  unsigned(0 downto 0);
o1 : out unsigned(0 downto 0);
o2 : out unsigned(0 downto 0);
o3 : out unsigned(71 downto 0));
end component cf_fft_256_18_18;
begin
n1 <= s27_1(6 downto 6) &
  s27_1(5 downto 5) &
  s27_1(4 downto 4) &
  s27_1(3 downto 3) &
  s27_1(2 downto 2) &
  s27_1(1 downto 1) &
  s27_1(0 downto 0);
n2 <= s25_1 & s25_2;
process (clock_c) begin
  if rising_edge(clock_c) then
    if i5 = "1" then
      n3 <= "0";
    elsif i4 = "1" then
      n3 <= s27_2;
    end if;
  end if;
end process;
process (clock_c) begin
  if rising_edge(clock_c) then
    if i5 = "1" then
      n4 <= "0";
    elsif i4 = "1" then
      n4 <= n3;
    end if;
  end if;
end process;
process (clock_c) begin
  if rising_edge(clock_c) then
    if i5 = "1" then
      n5 <= "0";
    elsif i4 = "1" then
      n5 <= n4;
    end if;
  end if;
end process;
process (clock_c) begin
  if rising_edge(clock_c) then
    if i5 = "1" then
      n6 <= "0";
    elsif i4 = "1" then
      n6 <= n5;
    end if;
  end if;
end process;
n7 <= s27_1(6 downto 6) &
  s27_1(5 downto 5) &
  s27_1(4 downto 4) &
  s27_1(3 downto 3) &
  s27_1(2 downto 2) &
  s27_1(1 downto 1);
process (clock_c) begin
  if rising_edge(clock_c) then
    if i5 = "1" then
      n8 <= "000000";
    elsif i4 = "1" then
      n8 <= n7;
    end if;
  end if;
end process;
process (clock_c) begin
  if rising_edge(clock_c) then
    if i5 = "1" then
      n9 <= "000000";
    elsif i4 = "1" then
      n9 <= n8;
    end if;
  end if;
end process;
process (clock_c) begin
  if rising_edge(clock_c) then
    if i5 = "1" then
      n10 <= "000000";
    elsif i4 = "1" then
      n10 <= n9;
    end if;
  end if;
end process;
process (clock_c) begin
  if rising_edge(clock_c) then
    if i5 = "1" then
      n11 <= "000000";
    elsif i4 = "1" then
      n11 <= n10;
    end if;
  end if;
end process;
n12 <= s27_1(0 downto 0);
process (clock_c) begin
  if rising_edge(clock_c) then
    if i5 = "1" then
      n13 <= "0";
    elsif i4 = "1" then
      n13 <= n12;
    end if;
  end if;
end process;
process (clock_c) begin
  if rising_edge(clock_c) then
    if i5 = "1" then
      n14 <= "0";
    elsif i4 = "1" then
      n14 <= n13;
    end if;
  end if;
end process;
process (clock_c) begin
  if rising_edge(clock_c) then
    if i5 = "1" then
      n15 <= "0";
    elsif i4 = "1" then
      n15 <= n14;
    end if;
  end if;
end process;
process (clock_c) begin
  if rising_edge(clock_c) then
    if i5 = "1" then
      n16 <= "0";
    elsif i4 = "1" then
      n16 <= n15;
    end if;
  end if;
end process;
n17 <= not n16;
n18 <= s29_2 & s29_1;
n19 <= s29_3(71 downto 71) &
  s29_3(70 downto 70) &
  s29_3(69 downto 69) &
  s29_3(68 downto 68) &
  s29_3(67 downto 67) &
  s29_3(66 downto 66) &
  s29_3(65 downto 65) &
  s29_3(64 downto 64) &
  s29_3(63 downto 63) &
  s29_3(62 downto 62) &
  s29_3(61 downto 61) &
  s29_3(60 downto 60) &
  s29_3(59 downto 59) &
  s29_3(58 downto 58) &
  s29_3(57 downto 57) &
  s29_3(56 downto 56) &
  s29_3(55 downto 55) &
  s29_3(54 downto 54) &
  s29_3(53 downto 53) &
  s29_3(52 downto 52) &
  s29_3(51 downto 51) &
  s29_3(50 downto 50) &
  s29_3(49 downto 49) &
  s29_3(48 downto 48) &
  s29_3(47 downto 47) &
  s29_3(46 downto 46) &
  s29_3(45 downto 45) &
  s29_3(44 downto 44) &
  s29_3(43 downto 43) &
  s29_3(42 downto 42) &
  s29_3(41 downto 41) &
  s29_3(40 downto 40) &
  s29_3(39 downto 39) &
  s29_3(38 downto 38) &
  s29_3(37 downto 37) &
  s29_3(36 downto 36);
n20 <= s29_3(35 downto 35) &
  s29_3(34 downto 34) &
  s29_3(33 downto 33) &
  s29_3(32 downto 32) &
  s29_3(31 downto 31) &
  s29_3(30 downto 30) &
  s29_3(29 downto 29) &
  s29_3(28 downto 28) &
  s29_3(27 downto 27) &
  s29_3(26 downto 26) &
  s29_3(25 downto 25) &
  s29_3(24 downto 24) &
  s29_3(23 downto 23) &
  s29_3(22 downto 22) &
  s29_3(21 downto 21) &
  s29_3(20 downto 20) &
  s29_3(19 downto 19) &
  s29_3(18 downto 18) &
  s29_3(17 downto 17) &
  s29_3(16 downto 16) &
  s29_3(15 downto 15) &
  s29_3(14 downto 14) &
  s29_3(13 downto 13) &
  s29_3(12 downto 12) &
  s29_3(11 downto 11) &
  s29_3(10 downto 10) &
  s29_3(9 downto 9) &
  s29_3(8 downto 8) &
  s29_3(7 downto 7) &
  s29_3(6 downto 6) &
  s29_3(5 downto 5) &
  s29_3(4 downto 4) &
  s29_3(3 downto 3) &
  s29_3(2 downto 2) &
  s29_3(1 downto 1) &
  s29_3(0 downto 0);
n21 <= s28_1(71 downto 71) &
  s28_1(70 downto 70) &
  s28_1(69 downto 69) &
  s28_1(68 downto 68) &
  s28_1(67 downto 67) &
  s28_1(66 downto 66) &
  s28_1(65 downto 65) &
  s28_1(64 downto 64) &
  s28_1(63 downto 63) &
  s28_1(62 downto 62) &
  s28_1(61 downto 61) &
  s28_1(60 downto 60) &
  s28_1(59 downto 59) &
  s28_1(58 downto 58) &
  s28_1(57 downto 57) &
  s28_1(56 downto 56) &
  s28_1(55 downto 55) &
  s28_1(54 downto 54) &
  s28_1(53 downto 53) &
  s28_1(52 downto 52) &
  s28_1(51 downto 51) &
  s28_1(50 downto 50) &
  s28_1(49 downto 49) &
  s28_1(48 downto 48) &
  s28_1(47 downto 47) &
  s28_1(46 downto 46) &
  s28_1(45 downto 45) &
  s28_1(44 downto 44) &
  s28_1(43 downto 43) &
  s28_1(42 downto 42) &
  s28_1(41 downto 41) &
  s28_1(40 downto 40) &
  s28_1(39 downto 39) &
  s28_1(38 downto 38) &
  s28_1(37 downto 37) &
  s28_1(36 downto 36);
n22 <= s28_1(35 downto 35) &
  s28_1(34 downto 34) &
  s28_1(33 downto 33) &
  s28_1(32 downto 32) &
  s28_1(31 downto 31) &
  s28_1(30 downto 30) &
  s28_1(29 downto 29) &
  s28_1(28 downto 28) &
  s28_1(27 downto 27) &
  s28_1(26 downto 26) &
  s28_1(25 downto 25) &
  s28_1(24 downto 24) &
  s28_1(23 downto 23) &
  s28_1(22 downto 22) &
  s28_1(21 downto 21) &
  s28_1(20 downto 20) &
  s28_1(19 downto 19) &
  s28_1(18 downto 18) &
  s28_1(17 downto 17) &
  s28_1(16 downto 16) &
  s28_1(15 downto 15) &
  s28_1(14 downto 14) &
  s28_1(13 downto 13) &
  s28_1(12 downto 12) &
  s28_1(11 downto 11) &
  s28_1(10 downto 10) &
  s28_1(9 downto 9) &
  s28_1(8 downto 8) &
  s28_1(7 downto 7) &
  s28_1(6 downto 6) &
  s28_1(5 downto 5) &
  s28_1(4 downto 4) &
  s28_1(3 downto 3) &
  s28_1(2 downto 2) &
  s28_1(1 downto 1) &
  s28_1(0 downto 0);
n23 <= n20 when s26_1 = "1" else n19;
n24 <= n22 when s26_1 = "1" else n21;
s25 : cf_fft_256_18_15 port map (clock_c, i2, i3, n1, i4, i5, s25_1, s25_2);
s26 : cf_fft_256_18_30 port map (clock_c, n18, i4, i5, s26_1);
s27 : cf_fft_256_18_21 port map (clock_c, i1, i4, i5, s27_1, s27_2);
s28 : cf_fft_256_18_17 port map (clock_c, n2, n6, n11, n16, i4, i5, s28_1);
s29 : cf_fft_256_18_18 port map (clock_c, n2, n6, n11, n17, i4, i5, s29_1, s29_2, s29_3);
o3 <= n24;
o2 <= n23;
o1 <= s29_1;
end architecture rtl;

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
entity cf_fft_256_18_13 is
port (
clock_c : in std_logic;
i1 : in  unsigned(35 downto 0);
i2 : in  unsigned(35 downto 0);
i3 : in  unsigned(4 downto 0);
i4 : in  unsigned(0 downto 0);
i5 : in  unsigned(0 downto 0);
o1 : out unsigned(35 downto 0);
o2 : out unsigned(35 downto 0));
end entity cf_fft_256_18_13;
architecture rtl of cf_fft_256_18_13 is
signal n1 : unsigned(35 downto 0) := "000000000000000000000000000000000000";
signal n2 : unsigned(17 downto 0);
signal n3 : unsigned(17 downto 0);
signal n4 : unsigned(35 downto 0) := "000000000000000000000000000000000000";
signal n5 : unsigned(17 downto 0);
signal n6 : unsigned(17 downto 0);
signal n7 : unsigned(17 downto 0) := "000000000000000000";
signal n8 : unsigned(17 downto 0) := "000000000000000000";
signal n9 : unsigned(17 downto 0) := "000000000000000000";
signal n10 : unsigned(17 downto 0) := "000000000000000000";
signal n11 : unsigned(35 downto 0) := "000000000000000000000000000000000000";
signal n12 : unsigned(17 downto 0);
signal n13 : unsigned(17 downto 0);
signal n14 : unsigned(35 downto 0);
signal n15 : unsigned(17 downto 0);
signal n16 : unsigned(17 downto 0) := "000000000000000000";
signal n17 : unsigned(35 downto 0);
signal n18 : unsigned(17 downto 0);
signal n19 : unsigned(17 downto 0) := "000000000000000000";
signal n20 : unsigned(17 downto 0);
signal n21 : unsigned(17 downto 0) := "000000000000000000";
signal n22 : unsigned(35 downto 0);
signal n23 : unsigned(17 downto 0);
signal n24 : unsigned(17 downto 0) := "000000000000000000";
signal n25 : unsigned(35 downto 0);
signal n26 : unsigned(17 downto 0);
signal n27 : unsigned(17 downto 0) := "000000000000000000";
signal n28 : unsigned(17 downto 0);
signal n29 : unsigned(17 downto 0) := "000000000000000000";
signal n30 : unsigned(17 downto 0);
signal n31 : unsigned(17 downto 0);
signal n32 : unsigned(35 downto 0);
signal n33 : unsigned(35 downto 0) := "000000000000000000000000000000000000";
signal n34 : unsigned(17 downto 0);
signal n35 : unsigned(17 downto 0);
signal n36 : unsigned(35 downto 0);
signal n37 : unsigned(35 downto 0) := "000000000000000000000000000000000000";
begin
process (clock_c) begin
  if rising_edge(clock_c) then
    if i5 = "1" then
      n1 <= "000000000000000000000000000000000000";
    elsif i4 = "1" then
      n1 <= i1;
    end if;
  end if;
end process;
n2 <= n1(35 downto 35) &
  n1(34 downto 34) &
  n1(33 downto 33) &
  n1(32 downto 32) &
  n1(31 downto 31) &
  n1(30 downto 30) &
  n1(29 downto 29) &
  n1(28 downto 28) &
  n1(27 downto 27) &
  n1(26 downto 26) &
  n1(25 downto 25) &
  n1(24 downto 24) &
  n1(23 downto 23) &
  n1(22 downto 22) &
  n1(21 downto 21) &
  n1(20 downto 20) &
  n1(19 downto 19) &
  n1(18 downto 18);
n3 <= n1(17 downto 17) &
  n1(16 downto 16) &
  n1(15 downto 15) &
  n1(14 downto 14) &
  n1(13 downto 13) &
  n1(12 downto 12) &
  n1(11 downto 11) &
  n1(10 downto 10) &
  n1(9 downto 9) &
  n1(8 downto 8) &
  n1(7 downto 7) &
  n1(6 downto 6) &
  n1(5 downto 5) &
  n1(4 downto 4) &
  n1(3 downto 3) &
  n1(2 downto 2) &
  n1(1 downto 1) &
  n1(0 downto 0);
process (clock_c) begin
  if rising_edge(clock_c) then
    if i5 = "1" then
      n4 <= "000000000000000000000000000000000000";
    elsif i4 = "1" then
      n4 <= i2;
    end if;
  end if;
end process;
n5 <= n4(35 downto 35) &
  n4(34 downto 34) &
  n4(33 downto 33) &
  n4(32 downto 32) &
  n4(31 downto 31) &
  n4(30 downto 30) &
  n4(29 downto 29) &
  n4(28 downto 28) &
  n4(27 downto 27) &
  n4(26 downto 26) &
  n4(25 downto 25) &
  n4(24 downto 24) &
  n4(23 downto 23) &
  n4(22 downto 22) &
  n4(21 downto 21) &
  n4(20 downto 20) &
  n4(19 downto 19) &
  n4(18 downto 18);
n6 <= n4(17 downto 17) &
  n4(16 downto 16) &
  n4(15 downto 15) &
  n4(14 downto 14) &
  n4(13 downto 13) &
  n4(12 downto 12) &
  n4(11 downto 11) &
  n4(10 downto 10) &
  n4(9 downto 9) &
  n4(8 downto 8) &
  n4(7 downto 7) &
  n4(6 downto 6) &
  n4(5 downto 5) &
  n4(4 downto 4) &
  n4(3 downto 3) &
  n4(2 downto 2) &
  n4(1 downto 1) &
  n4(0 downto 0);
process (clock_c) begin
  if rising_edge(clock_c) then
    if i5 = "1" then
      n7 <= "000000000000000000";
    elsif i4 = "1" then
      n7 <= n2;
    end if;
  end if;
end process;
process (clock_c) begin
  if rising_edge(clock_c) then
    if i5 = "1" then
      n8 <= "000000000000000000";
    elsif i4 = "1" then
      n8 <= n7;
    end if;
  end if;
end process;
process (clock_c) begin
  if rising_edge(clock_c) then
    if i5 = "1" then
      n9 <= "000000000000000000";
    elsif i4 = "1" then
      n9 <= n3;
    end if;
  end if;
end process;
process (clock_c) begin
  if rising_edge(clock_c) then
    if i5 = "1" then
      n10 <= "000000000000000000";
    elsif i4 = "1" then
      n10 <= n9;
    end if;
  end if;
end process;
process (clock_c) begin
  if rising_edge(clock_c) then 
    if i4 = "1" then
      case i3 is
        when "00000" => n11 <= "011111111111111111000000000000000000";
        when "00001" => n11 <= "011111110110001000111100110111010000";
        when "00010" => n11 <= "011111011000101001111001110000011101";
        when "00011" => n11 <= "011110100111110100110110101101011111";
        when "00100" => n11 <= "011101100100000110110011110000010000";
        when "00101" => n11 <= "011100001110001011110000111010100101";
        when "00110" => n11 <= "011010100110110110101110001110001100";
        when "00111" => n11 <= "011000101111001000101011101100110000";
        when "01000" => n11 <= "010110101000001001101001010111110110";
        when "01001" => n11 <= "010100010011001111100111010000110111";
        when "01010" => n11 <= "010001110001110011100101011001001001";
        when "01011" => n11 <= "001111000101011010100011110001110100";
        when "01100" => n11 <= "001100001111101111100010011011111001";
        when "01101" => n11 <= "001001010010100000100001011000001011";
        when "01110" => n11 <= "000110001111100010100000100111010110";
        when "01111" => n11 <= "000011001000101111100000001001110111";
        when "10000" => n11 <= "000000000000000000100000000000000000";
        when "10001" => n11 <= "111100110111010000100000001001110111";
        when "10010" => n11 <= "111001110000011101100000100111010110";
        when "10011" => n11 <= "110110101101011111100001011000001011";
        when "10100" => n11 <= "110011110000010000100010011011111001";
        when "10101" => n11 <= "110000111010100101100011110001110100";
        when "10110" => n11 <= "101110001110001100100101011001001001";
        when "10111" => n11 <= "101011101100110000100111010000110111";
        when "11000" => n11 <= "101001010111110110101001010111110110";
        when "11001" => n11 <= "100111010000110111101011101100110000";
        when "11010" => n11 <= "100101011001001001101110001110001100";
        when "11011" => n11 <= "100011110001110100110000111010100101";
        when "11100" => n11 <= "100010011011111001110011110000010000";
        when "11101" => n11 <= "100001011000001011110110101101011111";
        when "11110" => n11 <= "100000100111010110111001110000011101";
        when "11111" => n11 <= "100000001001110111111100110111010000";
        when others => n11 <= "XXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX";
      end case;
    end if;
  end if;
end process;
n12 <= n11(35 downto 35) &
  n11(34 downto 34) &
  n11(33 downto 33) &
  n11(32 downto 32) &
  n11(31 downto 31) &
  n11(30 downto 30) &
  n11(29 downto 29) &
  n11(28 downto 28) &
  n11(27 downto 27) &
  n11(26 downto 26) &
  n11(25 downto 25) &
  n11(24 downto 24) &
  n11(23 downto 23) &
  n11(22 downto 22) &
  n11(21 downto 21) &
  n11(20 downto 20) &
  n11(19 downto 19) &
  n11(18 downto 18);
n13 <= n11(17 downto 17) &
  n11(16 downto 16) &
  n11(15 downto 15) &
  n11(14 downto 14) &
  n11(13 downto 13) &
  n11(12 downto 12) &
  n11(11 downto 11) &
  n11(10 downto 10) &
  n11(9 downto 9) &
  n11(8 downto 8) &
  n11(7 downto 7) &
  n11(6 downto 6) &
  n11(5 downto 5) &
  n11(4 downto 4) &
  n11(3 downto 3) &
  n11(2 downto 2) &
  n11(1 downto 1) &
  n11(0 downto 0);
n14 <= unsigned(signed(n5) * signed(n12));
n15 <= n14(34 downto 34) &
  n14(33 downto 33) &
  n14(32 downto 32) &
  n14(31 downto 31) &
  n14(30 downto 30) &
  n14(29 downto 29) &
  n14(28 downto 28) &
  n14(27 downto 27) &
  n14(26 downto 26) &
  n14(25 downto 25) &
  n14(24 downto 24) &
  n14(23 downto 23) &
  n14(22 downto 22) &
  n14(21 downto 21) &
  n14(20 downto 20) &
  n14(19 downto 19) &
  n14(18 downto 18) &
  n14(17 downto 17);
process (clock_c) begin
  if rising_edge(clock_c) then
    if i5 = "1" then
      n16 <= "000000000000000000";
    elsif i4 = "1" then
      n16 <= n15;
    end if;
  end if;
end process;
n17 <= unsigned(signed(n6) * signed(n13));
n18 <= n17(34 downto 34) &
  n17(33 downto 33) &
  n17(32 downto 32) &
  n17(31 downto 31) &
  n17(30 downto 30) &
  n17(29 downto 29) &
  n17(28 downto 28) &
  n17(27 downto 27) &
  n17(26 downto 26) &
  n17(25 downto 25) &
  n17(24 downto 24) &
  n17(23 downto 23) &
  n17(22 downto 22) &
  n17(21 downto 21) &
  n17(20 downto 20) &
  n17(19 downto 19) &
  n17(18 downto 18) &
  n17(17 downto 17);
process (clock_c) begin
  if rising_edge(clock_c) then
    if i5 = "1" then
      n19 <= "000000000000000000";
    elsif i4 = "1" then
      n19 <= n18;
    end if;
  end if;
end process;
n20 <= n16 - n19;
process (clock_c) begin
  if rising_edge(clock_c) then
    if i5 = "1" then
      n21 <= "000000000000000000";
    elsif i4 = "1" then
      n21 <= n20;
    end if;
  end if;
end process;
n22 <= unsigned(signed(n5) * signed(n13));
n23 <= n22(34 downto 34) &
  n22(33 downto 33) &
  n22(32 downto 32) &
  n22(31 downto 31) &
  n22(30 downto 30) &
  n22(29 downto 29) &
  n22(28 downto 28) &
  n22(27 downto 27) &
  n22(26 downto 26) &
  n22(25 downto 25) &
  n22(24 downto 24) &
  n22(23 downto 23) &
  n22(22 downto 22) &
  n22(21 downto 21) &
  n22(20 downto 20) &
  n22(19 downto 19) &
  n22(18 downto 18) &
  n22(17 downto 17);
process (clock_c) begin
  if rising_edge(clock_c) then
    if i5 = "1" then
      n24 <= "000000000000000000";
    elsif i4 = "1" then
      n24 <= n23;
    end if;
  end if;
end process;
n25 <= unsigned(signed(n6) * signed(n12));
n26 <= n25(34 downto 34) &
  n25(33 downto 33) &
  n25(32 downto 32) &
  n25(31 downto 31) &
  n25(30 downto 30) &
  n25(29 downto 29) &
  n25(28 downto 28) &
  n25(27 downto 27) &
  n25(26 downto 26) &
  n25(25 downto 25) &
  n25(24 downto 24) &
  n25(23 downto 23) &
  n25(22 downto 22) &
  n25(21 downto 21) &
  n25(20 downto 20) &
  n25(19 downto 19) &
  n25(18 downto 18) &
  n25(17 downto 17);
process (clock_c) begin
  if rising_edge(clock_c) then
    if i5 = "1" then
      n27 <= "000000000000000000";
    elsif i4 = "1" then
      n27 <= n26;
    end if;
  end if;
end process;
n28 <= n24 + n27;
process (clock_c) begin
  if rising_edge(clock_c) then
    if i5 = "1" then
      n29 <= "000000000000000000";
    elsif i4 = "1" then
      n29 <= n28;
    end if;
  end if;
end process;
n30 <= n8 + n21;
n31 <= n10 + n29;
n32 <= n30 & n31;
process (clock_c) begin
  if rising_edge(clock_c) then
    if i5 = "1" then
      n33 <= "000000000000000000000000000000000000";
    elsif i4 = "1" then
      n33 <= n32;
    end if;
  end if;
end process;
n34 <= n8 - n21;
n35 <= n10 - n29;
n36 <= n34 & n35;
process (clock_c) begin
  if rising_edge(clock_c) then
    if i5 = "1" then
      n37 <= "000000000000000000000000000000000000";
    elsif i4 = "1" then
      n37 <= n36;
    end if;
  end if;
end process;
o2 <= n37;
o1 <= n33;
end architecture rtl;

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
entity cf_fft_256_18_12 is
port (
clock_c : in std_logic;
i1 : in  unsigned(0 downto 0);
i2 : in  unsigned(35 downto 0);
i3 : in  unsigned(35 downto 0);
i4 : in  unsigned(0 downto 0);
i5 : in  unsigned(0 downto 0);
o1 : out unsigned(0 downto 0);
o2 : out unsigned(35 downto 0);
o3 : out unsigned(35 downto 0));
end entity cf_fft_256_18_12;
architecture rtl of cf_fft_256_18_12 is
signal n1 : unsigned(4 downto 0);
signal n2 : unsigned(71 downto 0);
signal n3 : unsigned(0 downto 0) := "0";
signal n4 : unsigned(0 downto 0) := "0";
signal n5 : unsigned(0 downto 0) := "0";
signal n6 : unsigned(0 downto 0) := "0";
signal n7 : unsigned(5 downto 0);
signal n8 : unsigned(5 downto 0) := "000000";
signal n9 : unsigned(5 downto 0) := "000000";
signal n10 : unsigned(5 downto 0) := "000000";
signal n11 : unsigned(5 downto 0) := "000000";
signal n12 : unsigned(0 downto 0);
signal n13 : unsigned(0 downto 0) := "0";
signal n14 : unsigned(0 downto 0) := "0";
signal n15 : unsigned(0 downto 0) := "0";
signal n16 : unsigned(0 downto 0) := "0";
signal n17 : unsigned(0 downto 0);
signal n18 : unsigned(1 downto 0);
signal n19 : unsigned(35 downto 0);
signal n20 : unsigned(35 downto 0);
signal n21 : unsigned(35 downto 0);
signal n22 : unsigned(35 downto 0);
signal n23 : unsigned(35 downto 0);
signal n24 : unsigned(35 downto 0);
signal s25_1 : unsigned(0 downto 0);
signal s26_1 : unsigned(35 downto 0);
signal s26_2 : unsigned(35 downto 0);
signal s27_1 : unsigned(6 downto 0);
signal s27_2 : unsigned(0 downto 0);
signal s28_1 : unsigned(0 downto 0);
signal s28_2 : unsigned(0 downto 0);
signal s28_3 : unsigned(71 downto 0);
signal s29_1 : unsigned(71 downto 0);
component cf_fft_256_18_30 is
port (
clock_c : in std_logic;
i1 : in  unsigned(1 downto 0);
i2 : in  unsigned(0 downto 0);
i3 : in  unsigned(0 downto 0);
o1 : out unsigned(0 downto 0));
end component cf_fft_256_18_30;
component cf_fft_256_18_13 is
port (
clock_c : in std_logic;
i1 : in  unsigned(35 downto 0);
i2 : in  unsigned(35 downto 0);
i3 : in  unsigned(4 downto 0);
i4 : in  unsigned(0 downto 0);
i5 : in  unsigned(0 downto 0);
o1 : out unsigned(35 downto 0);
o2 : out unsigned(35 downto 0));
end component cf_fft_256_18_13;
component cf_fft_256_18_21 is
port (
clock_c : in std_logic;
i1 : in  unsigned(0 downto 0);
i2 : in  unsigned(0 downto 0);
i3 : in  unsigned(0 downto 0);
o1 : out unsigned(6 downto 0);
o2 : out unsigned(0 downto 0));
end component cf_fft_256_18_21;
component cf_fft_256_18_18 is
port (
clock_c : in std_logic;
i1 : in  unsigned(71 downto 0);
i2 : in  unsigned(0 downto 0);
i3 : in  unsigned(5 downto 0);
i4 : in  unsigned(0 downto 0);
i5 : in  unsigned(0 downto 0);
i6 : in  unsigned(0 downto 0);
o1 : out unsigned(0 downto 0);
o2 : out unsigned(0 downto 0);
o3 : out unsigned(71 downto 0));
end component cf_fft_256_18_18;
component cf_fft_256_18_17 is
port (
clock_c : in std_logic;
i1 : in  unsigned(71 downto 0);
i2 : in  unsigned(0 downto 0);
i3 : in  unsigned(5 downto 0);
i4 : in  unsigned(0 downto 0);
i5 : in  unsigned(0 downto 0);
i6 : in  unsigned(0 downto 0);
o1 : out unsigned(71 downto 0));
end component cf_fft_256_18_17;
begin
n1 <= s27_1(6 downto 6) &
  s27_1(5 downto 5) &
  s27_1(4 downto 4) &
  s27_1(3 downto 3) &
  s27_1(2 downto 2);
n2 <= s26_1 & s26_2;
process (clock_c) begin
  if rising_edge(clock_c) then
    if i5 = "1" then
      n3 <= "0";
    elsif i4 = "1" then
      n3 <= s27_2;
    end if;
  end if;
end process;
process (clock_c) begin
  if rising_edge(clock_c) then
    if i5 = "1" then
      n4 <= "0";
    elsif i4 = "1" then
      n4 <= n3;
    end if;
  end if;
end process;
process (clock_c) begin
  if rising_edge(clock_c) then
    if i5 = "1" then
      n5 <= "0";
    elsif i4 = "1" then
      n5 <= n4;
    end if;
  end if;
end process;
process (clock_c) begin
  if rising_edge(clock_c) then
    if i5 = "1" then
      n6 <= "0";
    elsif i4 = "1" then
      n6 <= n5;
    end if;
  end if;
end process;
n7 <= s27_1(6 downto 6) &
  s27_1(5 downto 5) &
  s27_1(4 downto 4) &
  s27_1(3 downto 3) &
  s27_1(2 downto 2) &
  s27_1(1 downto 1);
process (clock_c) begin
  if rising_edge(clock_c) then
    if i5 = "1" then
      n8 <= "000000";
    elsif i4 = "1" then
      n8 <= n7;
    end if;
  end if;
end process;
process (clock_c) begin
  if rising_edge(clock_c) then
    if i5 = "1" then
      n9 <= "000000";
    elsif i4 = "1" then
      n9 <= n8;
    end if;
  end if;
end process;
process (clock_c) begin
  if rising_edge(clock_c) then
    if i5 = "1" then
      n10 <= "000000";
    elsif i4 = "1" then
      n10 <= n9;
    end if;
  end if;
end process;
process (clock_c) begin
  if rising_edge(clock_c) then
    if i5 = "1" then
      n11 <= "000000";
    elsif i4 = "1" then
      n11 <= n10;
    end if;
  end if;
end process;
n12 <= s27_1(0 downto 0);
process (clock_c) begin
  if rising_edge(clock_c) then
    if i5 = "1" then
      n13 <= "0";
    elsif i4 = "1" then
      n13 <= n12;
    end if;
  end if;
end process;
process (clock_c) begin
  if rising_edge(clock_c) then
    if i5 = "1" then
      n14 <= "0";
    elsif i4 = "1" then
      n14 <= n13;
    end if;
  end if;
end process;
process (clock_c) begin
  if rising_edge(clock_c) then
    if i5 = "1" then
      n15 <= "0";
    elsif i4 = "1" then
      n15 <= n14;
    end if;
  end if;
end process;
process (clock_c) begin
  if rising_edge(clock_c) then
    if i5 = "1" then
      n16 <= "0";
    elsif i4 = "1" then
      n16 <= n15;
    end if;
  end if;
end process;
n17 <= not n16;
n18 <= s28_2 & s28_1;
n19 <= s28_3(71 downto 71) &
  s28_3(70 downto 70) &
  s28_3(69 downto 69) &
  s28_3(68 downto 68) &
  s28_3(67 downto 67) &
  s28_3(66 downto 66) &
  s28_3(65 downto 65) &
  s28_3(64 downto 64) &
  s28_3(63 downto 63) &
  s28_3(62 downto 62) &
  s28_3(61 downto 61) &
  s28_3(60 downto 60) &
  s28_3(59 downto 59) &
  s28_3(58 downto 58) &
  s28_3(57 downto 57) &
  s28_3(56 downto 56) &
  s28_3(55 downto 55) &
  s28_3(54 downto 54) &
  s28_3(53 downto 53) &
  s28_3(52 downto 52) &
  s28_3(51 downto 51) &
  s28_3(50 downto 50) &
  s28_3(49 downto 49) &
  s28_3(48 downto 48) &
  s28_3(47 downto 47) &
  s28_3(46 downto 46) &
  s28_3(45 downto 45) &
  s28_3(44 downto 44) &
  s28_3(43 downto 43) &
  s28_3(42 downto 42) &
  s28_3(41 downto 41) &
  s28_3(40 downto 40) &
  s28_3(39 downto 39) &
  s28_3(38 downto 38) &
  s28_3(37 downto 37) &
  s28_3(36 downto 36);
n20 <= s28_3(35 downto 35) &
  s28_3(34 downto 34) &
  s28_3(33 downto 33) &
  s28_3(32 downto 32) &
  s28_3(31 downto 31) &
  s28_3(30 downto 30) &
  s28_3(29 downto 29) &
  s28_3(28 downto 28) &
  s28_3(27 downto 27) &
  s28_3(26 downto 26) &
  s28_3(25 downto 25) &
  s28_3(24 downto 24) &
  s28_3(23 downto 23) &
  s28_3(22 downto 22) &
  s28_3(21 downto 21) &
  s28_3(20 downto 20) &
  s28_3(19 downto 19) &
  s28_3(18 downto 18) &
  s28_3(17 downto 17) &
  s28_3(16 downto 16) &
  s28_3(15 downto 15) &
  s28_3(14 downto 14) &
  s28_3(13 downto 13) &
  s28_3(12 downto 12) &
  s28_3(11 downto 11) &
  s28_3(10 downto 10) &
  s28_3(9 downto 9) &
  s28_3(8 downto 8) &
  s28_3(7 downto 7) &
  s28_3(6 downto 6) &
  s28_3(5 downto 5) &
  s28_3(4 downto 4) &
  s28_3(3 downto 3) &
  s28_3(2 downto 2) &
  s28_3(1 downto 1) &
  s28_3(0 downto 0);
n21 <= s29_1(71 downto 71) &
  s29_1(70 downto 70) &
  s29_1(69 downto 69) &
  s29_1(68 downto 68) &
  s29_1(67 downto 67) &
  s29_1(66 downto 66) &
  s29_1(65 downto 65) &
  s29_1(64 downto 64) &
  s29_1(63 downto 63) &
  s29_1(62 downto 62) &
  s29_1(61 downto 61) &
  s29_1(60 downto 60) &
  s29_1(59 downto 59) &
  s29_1(58 downto 58) &
  s29_1(57 downto 57) &
  s29_1(56 downto 56) &
  s29_1(55 downto 55) &
  s29_1(54 downto 54) &
  s29_1(53 downto 53) &
  s29_1(52 downto 52) &
  s29_1(51 downto 51) &
  s29_1(50 downto 50) &
  s29_1(49 downto 49) &
  s29_1(48 downto 48) &
  s29_1(47 downto 47) &
  s29_1(46 downto 46) &
  s29_1(45 downto 45) &
  s29_1(44 downto 44) &
  s29_1(43 downto 43) &
  s29_1(42 downto 42) &
  s29_1(41 downto 41) &
  s29_1(40 downto 40) &
  s29_1(39 downto 39) &
  s29_1(38 downto 38) &
  s29_1(37 downto 37) &
  s29_1(36 downto 36);
n22 <= s29_1(35 downto 35) &
  s29_1(34 downto 34) &
  s29_1(33 downto 33) &
  s29_1(32 downto 32) &
  s29_1(31 downto 31) &
  s29_1(30 downto 30) &
  s29_1(29 downto 29) &
  s29_1(28 downto 28) &
  s29_1(27 downto 27) &
  s29_1(26 downto 26) &
  s29_1(25 downto 25) &
  s29_1(24 downto 24) &
  s29_1(23 downto 23) &
  s29_1(22 downto 22) &
  s29_1(21 downto 21) &
  s29_1(20 downto 20) &
  s29_1(19 downto 19) &
  s29_1(18 downto 18) &
  s29_1(17 downto 17) &
  s29_1(16 downto 16) &
  s29_1(15 downto 15) &
  s29_1(14 downto 14) &
  s29_1(13 downto 13) &
  s29_1(12 downto 12) &
  s29_1(11 downto 11) &
  s29_1(10 downto 10) &
  s29_1(9 downto 9) &
  s29_1(8 downto 8) &
  s29_1(7 downto 7) &
  s29_1(6 downto 6) &
  s29_1(5 downto 5) &
  s29_1(4 downto 4) &
  s29_1(3 downto 3) &
  s29_1(2 downto 2) &
  s29_1(1 downto 1) &
  s29_1(0 downto 0);
n23 <= n20 when s25_1 = "1" else n19;
n24 <= n22 when s25_1 = "1" else n21;
s25 : cf_fft_256_18_30 port map (clock_c, n18, i4, i5, s25_1);
s26 : cf_fft_256_18_13 port map (clock_c, i2, i3, n1, i4, i5, s26_1, s26_2);
s27 : cf_fft_256_18_21 port map (clock_c, i1, i4, i5, s27_1, s27_2);
s28 : cf_fft_256_18_18 port map (clock_c, n2, n6, n11, n17, i4, i5, s28_1, s28_2, s28_3);
s29 : cf_fft_256_18_17 port map (clock_c, n2, n6, n11, n16, i4, i5, s29_1);
o3 <= n24;
o2 <= n23;
o1 <= s28_1;
end architecture rtl;

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
entity cf_fft_256_18_11 is
port (
clock_c : in std_logic;
i1 : in  unsigned(35 downto 0);
i2 : in  unsigned(35 downto 0);
i3 : in  unsigned(3 downto 0);
i4 : in  unsigned(0 downto 0);
i5 : in  unsigned(0 downto 0);
o1 : out unsigned(35 downto 0);
o2 : out unsigned(35 downto 0));
end entity cf_fft_256_18_11;
architecture rtl of cf_fft_256_18_11 is
signal n1 : unsigned(35 downto 0) := "000000000000000000000000000000000000";
signal n2 : unsigned(17 downto 0);
signal n3 : unsigned(17 downto 0);
signal n4 : unsigned(35 downto 0) := "000000000000000000000000000000000000";
signal n5 : unsigned(17 downto 0);
signal n6 : unsigned(17 downto 0);
signal n7 : unsigned(17 downto 0) := "000000000000000000";
signal n8 : unsigned(17 downto 0) := "000000000000000000";
signal n9 : unsigned(17 downto 0) := "000000000000000000";
signal n10 : unsigned(17 downto 0) := "000000000000000000";
signal n11 : unsigned(35 downto 0) := "000000000000000000000000000000000000";
signal n12 : unsigned(17 downto 0);
signal n13 : unsigned(17 downto 0);
signal n14 : unsigned(35 downto 0);
signal n15 : unsigned(17 downto 0);
signal n16 : unsigned(17 downto 0) := "000000000000000000";
signal n17 : unsigned(35 downto 0);
signal n18 : unsigned(17 downto 0);
signal n19 : unsigned(17 downto 0) := "000000000000000000";
signal n20 : unsigned(17 downto 0);
signal n21 : unsigned(17 downto 0) := "000000000000000000";
signal n22 : unsigned(35 downto 0);
signal n23 : unsigned(17 downto 0);
signal n24 : unsigned(17 downto 0) := "000000000000000000";
signal n25 : unsigned(35 downto 0);
signal n26 : unsigned(17 downto 0);
signal n27 : unsigned(17 downto 0) := "000000000000000000";
signal n28 : unsigned(17 downto 0);
signal n29 : unsigned(17 downto 0) := "000000000000000000";
signal n30 : unsigned(17 downto 0);
signal n31 : unsigned(17 downto 0);
signal n32 : unsigned(35 downto 0);
signal n33 : unsigned(35 downto 0) := "000000000000000000000000000000000000";
signal n34 : unsigned(17 downto 0);
signal n35 : unsigned(17 downto 0);
signal n36 : unsigned(35 downto 0);
signal n37 : unsigned(35 downto 0) := "000000000000000000000000000000000000";
begin
process (clock_c) begin
  if rising_edge(clock_c) then
    if i5 = "1" then
      n1 <= "000000000000000000000000000000000000";
    elsif i4 = "1" then
      n1 <= i1;
    end if;
  end if;
end process;
n2 <= n1(35 downto 35) &
  n1(34 downto 34) &
  n1(33 downto 33) &
  n1(32 downto 32) &
  n1(31 downto 31) &
  n1(30 downto 30) &
  n1(29 downto 29) &
  n1(28 downto 28) &
  n1(27 downto 27) &
  n1(26 downto 26) &
  n1(25 downto 25) &
  n1(24 downto 24) &
  n1(23 downto 23) &
  n1(22 downto 22) &
  n1(21 downto 21) &
  n1(20 downto 20) &
  n1(19 downto 19) &
  n1(18 downto 18);
n3 <= n1(17 downto 17) &
  n1(16 downto 16) &
  n1(15 downto 15) &
  n1(14 downto 14) &
  n1(13 downto 13) &
  n1(12 downto 12) &
  n1(11 downto 11) &
  n1(10 downto 10) &
  n1(9 downto 9) &
  n1(8 downto 8) &
  n1(7 downto 7) &
  n1(6 downto 6) &
  n1(5 downto 5) &
  n1(4 downto 4) &
  n1(3 downto 3) &
  n1(2 downto 2) &
  n1(1 downto 1) &
  n1(0 downto 0);
process (clock_c) begin
  if rising_edge(clock_c) then
    if i5 = "1" then
      n4 <= "000000000000000000000000000000000000";
    elsif i4 = "1" then
      n4 <= i2;
    end if;
  end if;
end process;
n5 <= n4(35 downto 35) &
  n4(34 downto 34) &
  n4(33 downto 33) &
  n4(32 downto 32) &
  n4(31 downto 31) &
  n4(30 downto 30) &
  n4(29 downto 29) &
  n4(28 downto 28) &
  n4(27 downto 27) &
  n4(26 downto 26) &
  n4(25 downto 25) &
  n4(24 downto 24) &
  n4(23 downto 23) &
  n4(22 downto 22) &
  n4(21 downto 21) &
  n4(20 downto 20) &
  n4(19 downto 19) &
  n4(18 downto 18);
n6 <= n4(17 downto 17) &
  n4(16 downto 16) &
  n4(15 downto 15) &
  n4(14 downto 14) &
  n4(13 downto 13) &
  n4(12 downto 12) &
  n4(11 downto 11) &
  n4(10 downto 10) &
  n4(9 downto 9) &
  n4(8 downto 8) &
  n4(7 downto 7) &
  n4(6 downto 6) &
  n4(5 downto 5) &
  n4(4 downto 4) &
  n4(3 downto 3) &
  n4(2 downto 2) &
  n4(1 downto 1) &
  n4(0 downto 0);
process (clock_c) begin
  if rising_edge(clock_c) then
    if i5 = "1" then
      n7 <= "000000000000000000";
    elsif i4 = "1" then
      n7 <= n2;
    end if;
  end if;
end process;
process (clock_c) begin
  if rising_edge(clock_c) then
    if i5 = "1" then
      n8 <= "000000000000000000";
    elsif i4 = "1" then
      n8 <= n7;
    end if;
  end if;
end process;
process (clock_c) begin
  if rising_edge(clock_c) then
    if i5 = "1" then
      n9 <= "000000000000000000";
    elsif i4 = "1" then
      n9 <= n3;
    end if;
  end if;
end process;
process (clock_c) begin
  if rising_edge(clock_c) then
    if i5 = "1" then
      n10 <= "000000000000000000";
    elsif i4 = "1" then
      n10 <= n9;
    end if;
  end if;
end process;
process (clock_c) begin
  if rising_edge(clock_c) then 
    if i4 = "1" then
      case i3 is
        when "0000" => n11 <= "011111111111111111000000000000000000";
        when "0001" => n11 <= "011111011000101001111001110000011101";
        when "0010" => n11 <= "011101100100000110110011110000010000";
        when "0011" => n11 <= "011010100110110110101110001110001100";
        when "0100" => n11 <= "010110101000001001101001010111110110";
        when "0101" => n11 <= "010001110001110011100101011001001001";
        when "0110" => n11 <= "001100001111101111100010011011111001";
        when "0111" => n11 <= "000110001111100010100000100111010110";
        when "1000" => n11 <= "000000000000000000100000000000000000";
        when "1001" => n11 <= "111001110000011101100000100111010110";
        when "1010" => n11 <= "110011110000010000100010011011111001";
        when "1011" => n11 <= "101110001110001100100101011001001001";
        when "1100" => n11 <= "101001010111110110101001010111110110";
        when "1101" => n11 <= "100101011001001001101110001110001100";
        when "1110" => n11 <= "100010011011111001110011110000010000";
        when "1111" => n11 <= "100000100111010110111001110000011101";
        when others => n11 <= "XXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX";
      end case;
    end if;
  end if;
end process;
n12 <= n11(35 downto 35) &
  n11(34 downto 34) &
  n11(33 downto 33) &
  n11(32 downto 32) &
  n11(31 downto 31) &
  n11(30 downto 30) &
  n11(29 downto 29) &
  n11(28 downto 28) &
  n11(27 downto 27) &
  n11(26 downto 26) &
  n11(25 downto 25) &
  n11(24 downto 24) &
  n11(23 downto 23) &
  n11(22 downto 22) &
  n11(21 downto 21) &
  n11(20 downto 20) &
  n11(19 downto 19) &
  n11(18 downto 18);
n13 <= n11(17 downto 17) &
  n11(16 downto 16) &
  n11(15 downto 15) &
  n11(14 downto 14) &
  n11(13 downto 13) &
  n11(12 downto 12) &
  n11(11 downto 11) &
  n11(10 downto 10) &
  n11(9 downto 9) &
  n11(8 downto 8) &
  n11(7 downto 7) &
  n11(6 downto 6) &
  n11(5 downto 5) &
  n11(4 downto 4) &
  n11(3 downto 3) &
  n11(2 downto 2) &
  n11(1 downto 1) &
  n11(0 downto 0);
n14 <= unsigned(signed(n5) * signed(n12));
n15 <= n14(34 downto 34) &
  n14(33 downto 33) &
  n14(32 downto 32) &
  n14(31 downto 31) &
  n14(30 downto 30) &
  n14(29 downto 29) &
  n14(28 downto 28) &
  n14(27 downto 27) &
  n14(26 downto 26) &
  n14(25 downto 25) &
  n14(24 downto 24) &
  n14(23 downto 23) &
  n14(22 downto 22) &
  n14(21 downto 21) &
  n14(20 downto 20) &
  n14(19 downto 19) &
  n14(18 downto 18) &
  n14(17 downto 17);
process (clock_c) begin
  if rising_edge(clock_c) then
    if i5 = "1" then
      n16 <= "000000000000000000";
    elsif i4 = "1" then
      n16 <= n15;
    end if;
  end if;
end process;
n17 <= unsigned(signed(n6) * signed(n13));
n18 <= n17(34 downto 34) &
  n17(33 downto 33) &
  n17(32 downto 32) &
  n17(31 downto 31) &
  n17(30 downto 30) &
  n17(29 downto 29) &
  n17(28 downto 28) &
  n17(27 downto 27) &
  n17(26 downto 26) &
  n17(25 downto 25) &
  n17(24 downto 24) &
  n17(23 downto 23) &
  n17(22 downto 22) &
  n17(21 downto 21) &
  n17(20 downto 20) &
  n17(19 downto 19) &
  n17(18 downto 18) &
  n17(17 downto 17);
process (clock_c) begin
  if rising_edge(clock_c) then
    if i5 = "1" then
      n19 <= "000000000000000000";
    elsif i4 = "1" then
      n19 <= n18;
    end if;
  end if;
end process;
n20 <= n16 - n19;
process (clock_c) begin
  if rising_edge(clock_c) then
    if i5 = "1" then
      n21 <= "000000000000000000";
    elsif i4 = "1" then
      n21 <= n20;
    end if;
  end if;
end process;
n22 <= unsigned(signed(n5) * signed(n13));
n23 <= n22(34 downto 34) &
  n22(33 downto 33) &
  n22(32 downto 32) &
  n22(31 downto 31) &
  n22(30 downto 30) &
  n22(29 downto 29) &
  n22(28 downto 28) &
  n22(27 downto 27) &
  n22(26 downto 26) &
  n22(25 downto 25) &
  n22(24 downto 24) &
  n22(23 downto 23) &
  n22(22 downto 22) &
  n22(21 downto 21) &
  n22(20 downto 20) &
  n22(19 downto 19) &
  n22(18 downto 18) &
  n22(17 downto 17);
process (clock_c) begin
  if rising_edge(clock_c) then
    if i5 = "1" then
      n24 <= "000000000000000000";
    elsif i4 = "1" then
      n24 <= n23;
    end if;
  end if;
end process;
n25 <= unsigned(signed(n6) * signed(n12));
n26 <= n25(34 downto 34) &
  n25(33 downto 33) &
  n25(32 downto 32) &
  n25(31 downto 31) &
  n25(30 downto 30) &
  n25(29 downto 29) &
  n25(28 downto 28) &
  n25(27 downto 27) &
  n25(26 downto 26) &
  n25(25 downto 25) &
  n25(24 downto 24) &
  n25(23 downto 23) &
  n25(22 downto 22) &
  n25(21 downto 21) &
  n25(20 downto 20) &
  n25(19 downto 19) &
  n25(18 downto 18) &
  n25(17 downto 17);
process (clock_c) begin
  if rising_edge(clock_c) then
    if i5 = "1" then
      n27 <= "000000000000000000";
    elsif i4 = "1" then
      n27 <= n26;
    end if;
  end if;
end process;
n28 <= n24 + n27;
process (clock_c) begin
  if rising_edge(clock_c) then
    if i5 = "1" then
      n29 <= "000000000000000000";
    elsif i4 = "1" then
      n29 <= n28;
    end if;
  end if;
end process;
n30 <= n8 + n21;
n31 <= n10 + n29;
n32 <= n30 & n31;
process (clock_c) begin
  if rising_edge(clock_c) then
    if i5 = "1" then
      n33 <= "000000000000000000000000000000000000";
    elsif i4 = "1" then
      n33 <= n32;
    end if;
  end if;
end process;
n34 <= n8 - n21;
n35 <= n10 - n29;
n36 <= n34 & n35;
process (clock_c) begin
  if rising_edge(clock_c) then
    if i5 = "1" then
      n37 <= "000000000000000000000000000000000000";
    elsif i4 = "1" then
      n37 <= n36;
    end if;
  end if;
end process;
o2 <= n37;
o1 <= n33;
end architecture rtl;

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
entity cf_fft_256_18_10 is
port (
clock_c : in std_logic;
i1 : in  unsigned(0 downto 0);
i2 : in  unsigned(35 downto 0);
i3 : in  unsigned(35 downto 0);
i4 : in  unsigned(0 downto 0);
i5 : in  unsigned(0 downto 0);
o1 : out unsigned(0 downto 0);
o2 : out unsigned(35 downto 0);
o3 : out unsigned(35 downto 0));
end entity cf_fft_256_18_10;
architecture rtl of cf_fft_256_18_10 is
signal n1 : unsigned(3 downto 0);
signal n2 : unsigned(71 downto 0);
signal n3 : unsigned(0 downto 0) := "0";
signal n4 : unsigned(0 downto 0) := "0";
signal n5 : unsigned(0 downto 0) := "0";
signal n6 : unsigned(0 downto 0) := "0";
signal n7 : unsigned(5 downto 0);
signal n8 : unsigned(5 downto 0) := "000000";
signal n9 : unsigned(5 downto 0) := "000000";
signal n10 : unsigned(5 downto 0) := "000000";
signal n11 : unsigned(5 downto 0) := "000000";
signal n12 : unsigned(0 downto 0);
signal n13 : unsigned(0 downto 0) := "0";
signal n14 : unsigned(0 downto 0) := "0";
signal n15 : unsigned(0 downto 0) := "0";
signal n16 : unsigned(0 downto 0) := "0";
signal n17 : unsigned(0 downto 0);
signal n18 : unsigned(1 downto 0);
signal n19 : unsigned(35 downto 0);
signal n20 : unsigned(35 downto 0);
signal n21 : unsigned(35 downto 0);
signal n22 : unsigned(35 downto 0);
signal n23 : unsigned(35 downto 0);
signal n24 : unsigned(35 downto 0);
signal s25_1 : unsigned(0 downto 0);
signal s26_1 : unsigned(35 downto 0);
signal s26_2 : unsigned(35 downto 0);
signal s27_1 : unsigned(6 downto 0);
signal s27_2 : unsigned(0 downto 0);
signal s28_1 : unsigned(0 downto 0);
signal s28_2 : unsigned(0 downto 0);
signal s28_3 : unsigned(71 downto 0);
signal s29_1 : unsigned(71 downto 0);
component cf_fft_256_18_30 is
port (
clock_c : in std_logic;
i1 : in  unsigned(1 downto 0);
i2 : in  unsigned(0 downto 0);
i3 : in  unsigned(0 downto 0);
o1 : out unsigned(0 downto 0));
end component cf_fft_256_18_30;
component cf_fft_256_18_11 is
port (
clock_c : in std_logic;
i1 : in  unsigned(35 downto 0);
i2 : in  unsigned(35 downto 0);
i3 : in  unsigned(3 downto 0);
i4 : in  unsigned(0 downto 0);
i5 : in  unsigned(0 downto 0);
o1 : out unsigned(35 downto 0);
o2 : out unsigned(35 downto 0));
end component cf_fft_256_18_11;
component cf_fft_256_18_21 is
port (
clock_c : in std_logic;
i1 : in  unsigned(0 downto 0);
i2 : in  unsigned(0 downto 0);
i3 : in  unsigned(0 downto 0);
o1 : out unsigned(6 downto 0);
o2 : out unsigned(0 downto 0));
end component cf_fft_256_18_21;
component cf_fft_256_18_18 is
port (
clock_c : in std_logic;
i1 : in  unsigned(71 downto 0);
i2 : in  unsigned(0 downto 0);
i3 : in  unsigned(5 downto 0);
i4 : in  unsigned(0 downto 0);
i5 : in  unsigned(0 downto 0);
i6 : in  unsigned(0 downto 0);
o1 : out unsigned(0 downto 0);
o2 : out unsigned(0 downto 0);
o3 : out unsigned(71 downto 0));
end component cf_fft_256_18_18;
component cf_fft_256_18_17 is
port (
clock_c : in std_logic;
i1 : in  unsigned(71 downto 0);
i2 : in  unsigned(0 downto 0);
i3 : in  unsigned(5 downto 0);
i4 : in  unsigned(0 downto 0);
i5 : in  unsigned(0 downto 0);
i6 : in  unsigned(0 downto 0);
o1 : out unsigned(71 downto 0));
end component cf_fft_256_18_17;
begin
n1 <= s27_1(6 downto 6) &
  s27_1(5 downto 5) &
  s27_1(4 downto 4) &
  s27_1(3 downto 3);
n2 <= s26_1 & s26_2;
process (clock_c) begin
  if rising_edge(clock_c) then
    if i5 = "1" then
      n3 <= "0";
    elsif i4 = "1" then
      n3 <= s27_2;
    end if;
  end if;
end process;
process (clock_c) begin
  if rising_edge(clock_c) then
    if i5 = "1" then
      n4 <= "0";
    elsif i4 = "1" then
      n4 <= n3;
    end if;
  end if;
end process;
process (clock_c) begin
  if rising_edge(clock_c) then
    if i5 = "1" then
      n5 <= "0";
    elsif i4 = "1" then
      n5 <= n4;
    end if;
  end if;
end process;
process (clock_c) begin
  if rising_edge(clock_c) then
    if i5 = "1" then
      n6 <= "0";
    elsif i4 = "1" then
      n6 <= n5;
    end if;
  end if;
end process;
n7 <= s27_1(6 downto 6) &
  s27_1(5 downto 5) &
  s27_1(4 downto 4) &
  s27_1(3 downto 3) &
  s27_1(2 downto 2) &
  s27_1(1 downto 1);
process (clock_c) begin
  if rising_edge(clock_c) then
    if i5 = "1" then
      n8 <= "000000";
    elsif i4 = "1" then
      n8 <= n7;
    end if;
  end if;
end process;
process (clock_c) begin
  if rising_edge(clock_c) then
    if i5 = "1" then
      n9 <= "000000";
    elsif i4 = "1" then
      n9 <= n8;
    end if;
  end if;
end process;
process (clock_c) begin
  if rising_edge(clock_c) then
    if i5 = "1" then
      n10 <= "000000";
    elsif i4 = "1" then
      n10 <= n9;
    end if;
  end if;
end process;
process (clock_c) begin
  if rising_edge(clock_c) then
    if i5 = "1" then
      n11 <= "000000";
    elsif i4 = "1" then
      n11 <= n10;
    end if;
  end if;
end process;
n12 <= s27_1(0 downto 0);
process (clock_c) begin
  if rising_edge(clock_c) then
    if i5 = "1" then
      n13 <= "0";
    elsif i4 = "1" then
      n13 <= n12;
    end if;
  end if;
end process;
process (clock_c) begin
  if rising_edge(clock_c) then
    if i5 = "1" then
      n14 <= "0";
    elsif i4 = "1" then
      n14 <= n13;
    end if;
  end if;
end process;
process (clock_c) begin
  if rising_edge(clock_c) then
    if i5 = "1" then
      n15 <= "0";
    elsif i4 = "1" then
      n15 <= n14;
    end if;
  end if;
end process;
process (clock_c) begin
  if rising_edge(clock_c) then
    if i5 = "1" then
      n16 <= "0";
    elsif i4 = "1" then
      n16 <= n15;
    end if;
  end if;
end process;
n17 <= not n16;
n18 <= s28_2 & s28_1;
n19 <= s28_3(71 downto 71) &
  s28_3(70 downto 70) &
  s28_3(69 downto 69) &
  s28_3(68 downto 68) &
  s28_3(67 downto 67) &
  s28_3(66 downto 66) &
  s28_3(65 downto 65) &
  s28_3(64 downto 64) &
  s28_3(63 downto 63) &
  s28_3(62 downto 62) &
  s28_3(61 downto 61) &
  s28_3(60 downto 60) &
  s28_3(59 downto 59) &
  s28_3(58 downto 58) &
  s28_3(57 downto 57) &
  s28_3(56 downto 56) &
  s28_3(55 downto 55) &
  s28_3(54 downto 54) &
  s28_3(53 downto 53) &
  s28_3(52 downto 52) &
  s28_3(51 downto 51) &
  s28_3(50 downto 50) &
  s28_3(49 downto 49) &
  s28_3(48 downto 48) &
  s28_3(47 downto 47) &
  s28_3(46 downto 46) &
  s28_3(45 downto 45) &
  s28_3(44 downto 44) &
  s28_3(43 downto 43) &
  s28_3(42 downto 42) &
  s28_3(41 downto 41) &
  s28_3(40 downto 40) &
  s28_3(39 downto 39) &
  s28_3(38 downto 38) &
  s28_3(37 downto 37) &
  s28_3(36 downto 36);
n20 <= s28_3(35 downto 35) &
  s28_3(34 downto 34) &
  s28_3(33 downto 33) &
  s28_3(32 downto 32) &
  s28_3(31 downto 31) &
  s28_3(30 downto 30) &
  s28_3(29 downto 29) &
  s28_3(28 downto 28) &
  s28_3(27 downto 27) &
  s28_3(26 downto 26) &
  s28_3(25 downto 25) &
  s28_3(24 downto 24) &
  s28_3(23 downto 23) &
  s28_3(22 downto 22) &
  s28_3(21 downto 21) &
  s28_3(20 downto 20) &
  s28_3(19 downto 19) &
  s28_3(18 downto 18) &
  s28_3(17 downto 17) &
  s28_3(16 downto 16) &
  s28_3(15 downto 15) &
  s28_3(14 downto 14) &
  s28_3(13 downto 13) &
  s28_3(12 downto 12) &
  s28_3(11 downto 11) &
  s28_3(10 downto 10) &
  s28_3(9 downto 9) &
  s28_3(8 downto 8) &
  s28_3(7 downto 7) &
  s28_3(6 downto 6) &
  s28_3(5 downto 5) &
  s28_3(4 downto 4) &
  s28_3(3 downto 3) &
  s28_3(2 downto 2) &
  s28_3(1 downto 1) &
  s28_3(0 downto 0);
n21 <= s29_1(71 downto 71) &
  s29_1(70 downto 70) &
  s29_1(69 downto 69) &
  s29_1(68 downto 68) &
  s29_1(67 downto 67) &
  s29_1(66 downto 66) &
  s29_1(65 downto 65) &
  s29_1(64 downto 64) &
  s29_1(63 downto 63) &
  s29_1(62 downto 62) &
  s29_1(61 downto 61) &
  s29_1(60 downto 60) &
  s29_1(59 downto 59) &
  s29_1(58 downto 58) &
  s29_1(57 downto 57) &
  s29_1(56 downto 56) &
  s29_1(55 downto 55) &
  s29_1(54 downto 54) &
  s29_1(53 downto 53) &
  s29_1(52 downto 52) &
  s29_1(51 downto 51) &
  s29_1(50 downto 50) &
  s29_1(49 downto 49) &
  s29_1(48 downto 48) &
  s29_1(47 downto 47) &
  s29_1(46 downto 46) &
  s29_1(45 downto 45) &
  s29_1(44 downto 44) &
  s29_1(43 downto 43) &
  s29_1(42 downto 42) &
  s29_1(41 downto 41) &
  s29_1(40 downto 40) &
  s29_1(39 downto 39) &
  s29_1(38 downto 38) &
  s29_1(37 downto 37) &
  s29_1(36 downto 36);
n22 <= s29_1(35 downto 35) &
  s29_1(34 downto 34) &
  s29_1(33 downto 33) &
  s29_1(32 downto 32) &
  s29_1(31 downto 31) &
  s29_1(30 downto 30) &
  s29_1(29 downto 29) &
  s29_1(28 downto 28) &
  s29_1(27 downto 27) &
  s29_1(26 downto 26) &
  s29_1(25 downto 25) &
  s29_1(24 downto 24) &
  s29_1(23 downto 23) &
  s29_1(22 downto 22) &
  s29_1(21 downto 21) &
  s29_1(20 downto 20) &
  s29_1(19 downto 19) &
  s29_1(18 downto 18) &
  s29_1(17 downto 17) &
  s29_1(16 downto 16) &
  s29_1(15 downto 15) &
  s29_1(14 downto 14) &
  s29_1(13 downto 13) &
  s29_1(12 downto 12) &
  s29_1(11 downto 11) &
  s29_1(10 downto 10) &
  s29_1(9 downto 9) &
  s29_1(8 downto 8) &
  s29_1(7 downto 7) &
  s29_1(6 downto 6) &
  s29_1(5 downto 5) &
  s29_1(4 downto 4) &
  s29_1(3 downto 3) &
  s29_1(2 downto 2) &
  s29_1(1 downto 1) &
  s29_1(0 downto 0);
n23 <= n20 when s25_1 = "1" else n19;
n24 <= n22 when s25_1 = "1" else n21;
s25 : cf_fft_256_18_30 port map (clock_c, n18, i4, i5, s25_1);
s26 : cf_fft_256_18_11 port map (clock_c, i2, i3, n1, i4, i5, s26_1, s26_2);
s27 : cf_fft_256_18_21 port map (clock_c, i1, i4, i5, s27_1, s27_2);
s28 : cf_fft_256_18_18 port map (clock_c, n2, n6, n11, n17, i4, i5, s28_1, s28_2, s28_3);
s29 : cf_fft_256_18_17 port map (clock_c, n2, n6, n11, n16, i4, i5, s29_1);
o3 <= n24;
o2 <= n23;
o1 <= s28_1;
end architecture rtl;

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
entity cf_fft_256_18_9 is
port (
clock_c : in std_logic;
i1 : in  unsigned(35 downto 0);
i2 : in  unsigned(35 downto 0);
i3 : in  unsigned(2 downto 0);
i4 : in  unsigned(0 downto 0);
i5 : in  unsigned(0 downto 0);
o1 : out unsigned(35 downto 0);
o2 : out unsigned(35 downto 0));
end entity cf_fft_256_18_9;
architecture rtl of cf_fft_256_18_9 is
signal n1 : unsigned(35 downto 0) := "000000000000000000000000000000000000";
signal n2 : unsigned(17 downto 0);
signal n3 : unsigned(17 downto 0);
signal n4 : unsigned(35 downto 0) := "000000000000000000000000000000000000";
signal n5 : unsigned(17 downto 0);
signal n6 : unsigned(17 downto 0);
signal n7 : unsigned(17 downto 0) := "000000000000000000";
signal n8 : unsigned(17 downto 0) := "000000000000000000";
signal n9 : unsigned(17 downto 0) := "000000000000000000";
signal n10 : unsigned(17 downto 0) := "000000000000000000";
signal n11 : unsigned(35 downto 0) := "000000000000000000000000000000000000";
signal n12 : unsigned(17 downto 0);
signal n13 : unsigned(17 downto 0);
signal n14 : unsigned(35 downto 0);
signal n15 : unsigned(17 downto 0);
signal n16 : unsigned(17 downto 0) := "000000000000000000";
signal n17 : unsigned(35 downto 0);
signal n18 : unsigned(17 downto 0);
signal n19 : unsigned(17 downto 0) := "000000000000000000";
signal n20 : unsigned(17 downto 0);
signal n21 : unsigned(17 downto 0) := "000000000000000000";
signal n22 : unsigned(35 downto 0);
signal n23 : unsigned(17 downto 0);
signal n24 : unsigned(17 downto 0) := "000000000000000000";
signal n25 : unsigned(35 downto 0);
signal n26 : unsigned(17 downto 0);
signal n27 : unsigned(17 downto 0) := "000000000000000000";
signal n28 : unsigned(17 downto 0);
signal n29 : unsigned(17 downto 0) := "000000000000000000";
signal n30 : unsigned(17 downto 0);
signal n31 : unsigned(17 downto 0);
signal n32 : unsigned(35 downto 0);
signal n33 : unsigned(35 downto 0) := "000000000000000000000000000000000000";
signal n34 : unsigned(17 downto 0);
signal n35 : unsigned(17 downto 0);
signal n36 : unsigned(35 downto 0);
signal n37 : unsigned(35 downto 0) := "000000000000000000000000000000000000";
begin
process (clock_c) begin
  if rising_edge(clock_c) then
    if i5 = "1" then
      n1 <= "000000000000000000000000000000000000";
    elsif i4 = "1" then
      n1 <= i1;
    end if;
  end if;
end process;
n2 <= n1(35 downto 35) &
  n1(34 downto 34) &
  n1(33 downto 33) &
  n1(32 downto 32) &
  n1(31 downto 31) &
  n1(30 downto 30) &
  n1(29 downto 29) &
  n1(28 downto 28) &
  n1(27 downto 27) &
  n1(26 downto 26) &
  n1(25 downto 25) &
  n1(24 downto 24) &
  n1(23 downto 23) &
  n1(22 downto 22) &
  n1(21 downto 21) &
  n1(20 downto 20) &
  n1(19 downto 19) &
  n1(18 downto 18);
n3 <= n1(17 downto 17) &
  n1(16 downto 16) &
  n1(15 downto 15) &
  n1(14 downto 14) &
  n1(13 downto 13) &
  n1(12 downto 12) &
  n1(11 downto 11) &
  n1(10 downto 10) &
  n1(9 downto 9) &
  n1(8 downto 8) &
  n1(7 downto 7) &
  n1(6 downto 6) &
  n1(5 downto 5) &
  n1(4 downto 4) &
  n1(3 downto 3) &
  n1(2 downto 2) &
  n1(1 downto 1) &
  n1(0 downto 0);
process (clock_c) begin
  if rising_edge(clock_c) then
    if i5 = "1" then
      n4 <= "000000000000000000000000000000000000";
    elsif i4 = "1" then
      n4 <= i2;
    end if;
  end if;
end process;
n5 <= n4(35 downto 35) &
  n4(34 downto 34) &
  n4(33 downto 33) &
  n4(32 downto 32) &
  n4(31 downto 31) &
  n4(30 downto 30) &
  n4(29 downto 29) &
  n4(28 downto 28) &
  n4(27 downto 27) &
  n4(26 downto 26) &
  n4(25 downto 25) &
  n4(24 downto 24) &
  n4(23 downto 23) &
  n4(22 downto 22) &
  n4(21 downto 21) &
  n4(20 downto 20) &
  n4(19 downto 19) &
  n4(18 downto 18);
n6 <= n4(17 downto 17) &
  n4(16 downto 16) &
  n4(15 downto 15) &
  n4(14 downto 14) &
  n4(13 downto 13) &
  n4(12 downto 12) &
  n4(11 downto 11) &
  n4(10 downto 10) &
  n4(9 downto 9) &
  n4(8 downto 8) &
  n4(7 downto 7) &
  n4(6 downto 6) &
  n4(5 downto 5) &
  n4(4 downto 4) &
  n4(3 downto 3) &
  n4(2 downto 2) &
  n4(1 downto 1) &
  n4(0 downto 0);
process (clock_c) begin
  if rising_edge(clock_c) then
    if i5 = "1" then
      n7 <= "000000000000000000";
    elsif i4 = "1" then
      n7 <= n2;
    end if;
  end if;
end process;
process (clock_c) begin
  if rising_edge(clock_c) then
    if i5 = "1" then
      n8 <= "000000000000000000";
    elsif i4 = "1" then
      n8 <= n7;
    end if;
  end if;
end process;
process (clock_c) begin
  if rising_edge(clock_c) then
    if i5 = "1" then
      n9 <= "000000000000000000";
    elsif i4 = "1" then
      n9 <= n3;
    end if;
  end if;
end process;
process (clock_c) begin
  if rising_edge(clock_c) then
    if i5 = "1" then
      n10 <= "000000000000000000";
    elsif i4 = "1" then
      n10 <= n9;
    end if;
  end if;
end process;
process (clock_c) begin
  if rising_edge(clock_c) then 
    if i4 = "1" then
      case i3 is
        when "000" => n11 <= "011111111111111111000000000000000000";
        when "001" => n11 <= "011101100100000110110011110000010000";
        when "010" => n11 <= "010110101000001001101001010111110110";
        when "011" => n11 <= "001100001111101111100010011011111001";
        when "100" => n11 <= "000000000000000000100000000000000000";
        when "101" => n11 <= "110011110000010000100010011011111001";
        when "110" => n11 <= "101001010111110110101001010111110110";
        when "111" => n11 <= "100010011011111001110011110000010000";
        when others => n11 <= "XXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX";
      end case;
    end if;
  end if;
end process;
n12 <= n11(35 downto 35) &
  n11(34 downto 34) &
  n11(33 downto 33) &
  n11(32 downto 32) &
  n11(31 downto 31) &
  n11(30 downto 30) &
  n11(29 downto 29) &
  n11(28 downto 28) &
  n11(27 downto 27) &
  n11(26 downto 26) &
  n11(25 downto 25) &
  n11(24 downto 24) &
  n11(23 downto 23) &
  n11(22 downto 22) &
  n11(21 downto 21) &
  n11(20 downto 20) &
  n11(19 downto 19) &
  n11(18 downto 18);
n13 <= n11(17 downto 17) &
  n11(16 downto 16) &
  n11(15 downto 15) &
  n11(14 downto 14) &
  n11(13 downto 13) &
  n11(12 downto 12) &
  n11(11 downto 11) &
  n11(10 downto 10) &
  n11(9 downto 9) &
  n11(8 downto 8) &
  n11(7 downto 7) &
  n11(6 downto 6) &
  n11(5 downto 5) &
  n11(4 downto 4) &
  n11(3 downto 3) &
  n11(2 downto 2) &
  n11(1 downto 1) &
  n11(0 downto 0);
n14 <= unsigned(signed(n5) * signed(n12));
n15 <= n14(34 downto 34) &
  n14(33 downto 33) &
  n14(32 downto 32) &
  n14(31 downto 31) &
  n14(30 downto 30) &
  n14(29 downto 29) &
  n14(28 downto 28) &
  n14(27 downto 27) &
  n14(26 downto 26) &
  n14(25 downto 25) &
  n14(24 downto 24) &
  n14(23 downto 23) &
  n14(22 downto 22) &
  n14(21 downto 21) &
  n14(20 downto 20) &
  n14(19 downto 19) &
  n14(18 downto 18) &
  n14(17 downto 17);
process (clock_c) begin
  if rising_edge(clock_c) then
    if i5 = "1" then
      n16 <= "000000000000000000";
    elsif i4 = "1" then
      n16 <= n15;
    end if;
  end if;
end process;
n17 <= unsigned(signed(n6) * signed(n13));
n18 <= n17(34 downto 34) &
  n17(33 downto 33) &
  n17(32 downto 32) &
  n17(31 downto 31) &
  n17(30 downto 30) &
  n17(29 downto 29) &
  n17(28 downto 28) &
  n17(27 downto 27) &
  n17(26 downto 26) &
  n17(25 downto 25) &
  n17(24 downto 24) &
  n17(23 downto 23) &
  n17(22 downto 22) &
  n17(21 downto 21) &
  n17(20 downto 20) &
  n17(19 downto 19) &
  n17(18 downto 18) &
  n17(17 downto 17);
process (clock_c) begin
  if rising_edge(clock_c) then
    if i5 = "1" then
      n19 <= "000000000000000000";
    elsif i4 = "1" then
      n19 <= n18;
    end if;
  end if;
end process;
n20 <= n16 - n19;
process (clock_c) begin
  if rising_edge(clock_c) then
    if i5 = "1" then
      n21 <= "000000000000000000";
    elsif i4 = "1" then
      n21 <= n20;
    end if;
  end if;
end process;
n22 <= unsigned(signed(n5) * signed(n13));
n23 <= n22(34 downto 34) &
  n22(33 downto 33) &
  n22(32 downto 32) &
  n22(31 downto 31) &
  n22(30 downto 30) &
  n22(29 downto 29) &
  n22(28 downto 28) &
  n22(27 downto 27) &
  n22(26 downto 26) &
  n22(25 downto 25) &
  n22(24 downto 24) &
  n22(23 downto 23) &
  n22(22 downto 22) &
  n22(21 downto 21) &
  n22(20 downto 20) &
  n22(19 downto 19) &
  n22(18 downto 18) &
  n22(17 downto 17);
process (clock_c) begin
  if rising_edge(clock_c) then
    if i5 = "1" then
      n24 <= "000000000000000000";
    elsif i4 = "1" then
      n24 <= n23;
    end if;
  end if;
end process;
n25 <= unsigned(signed(n6) * signed(n12));
n26 <= n25(34 downto 34) &
  n25(33 downto 33) &
  n25(32 downto 32) &
  n25(31 downto 31) &
  n25(30 downto 30) &
  n25(29 downto 29) &
  n25(28 downto 28) &
  n25(27 downto 27) &
  n25(26 downto 26) &
  n25(25 downto 25) &
  n25(24 downto 24) &
  n25(23 downto 23) &
  n25(22 downto 22) &
  n25(21 downto 21) &
  n25(20 downto 20) &
  n25(19 downto 19) &
  n25(18 downto 18) &
  n25(17 downto 17);
process (clock_c) begin
  if rising_edge(clock_c) then
    if i5 = "1" then
      n27 <= "000000000000000000";
    elsif i4 = "1" then
      n27 <= n26;
    end if;
  end if;
end process;
n28 <= n24 + n27;
process (clock_c) begin
  if rising_edge(clock_c) then
    if i5 = "1" then
      n29 <= "000000000000000000";
    elsif i4 = "1" then
      n29 <= n28;
    end if;
  end if;
end process;
n30 <= n8 + n21;
n31 <= n10 + n29;
n32 <= n30 & n31;
process (clock_c) begin
  if rising_edge(clock_c) then
    if i5 = "1" then
      n33 <= "000000000000000000000000000000000000";
    elsif i4 = "1" then
      n33 <= n32;
    end if;
  end if;
end process;
n34 <= n8 - n21;
n35 <= n10 - n29;
n36 <= n34 & n35;
process (clock_c) begin
  if rising_edge(clock_c) then
    if i5 = "1" then
      n37 <= "000000000000000000000000000000000000";
    elsif i4 = "1" then
      n37 <= n36;
    end if;
  end if;
end process;
o2 <= n37;
o1 <= n33;
end architecture rtl;

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
entity cf_fft_256_18_8 is
port (
clock_c : in std_logic;
i1 : in  unsigned(0 downto 0);
i2 : in  unsigned(35 downto 0);
i3 : in  unsigned(35 downto 0);
i4 : in  unsigned(0 downto 0);
i5 : in  unsigned(0 downto 0);
o1 : out unsigned(0 downto 0);
o2 : out unsigned(35 downto 0);
o3 : out unsigned(35 downto 0));
end entity cf_fft_256_18_8;
architecture rtl of cf_fft_256_18_8 is
signal n1 : unsigned(2 downto 0);
signal n2 : unsigned(71 downto 0);
signal n3 : unsigned(0 downto 0) := "0";
signal n4 : unsigned(0 downto 0) := "0";
signal n5 : unsigned(0 downto 0) := "0";
signal n6 : unsigned(0 downto 0) := "0";
signal n7 : unsigned(5 downto 0);
signal n8 : unsigned(5 downto 0) := "000000";
signal n9 : unsigned(5 downto 0) := "000000";
signal n10 : unsigned(5 downto 0) := "000000";
signal n11 : unsigned(5 downto 0) := "000000";
signal n12 : unsigned(0 downto 0);
signal n13 : unsigned(0 downto 0) := "0";
signal n14 : unsigned(0 downto 0) := "0";
signal n15 : unsigned(0 downto 0) := "0";
signal n16 : unsigned(0 downto 0) := "0";
signal n17 : unsigned(0 downto 0);
signal n18 : unsigned(1 downto 0);
signal n19 : unsigned(35 downto 0);
signal n20 : unsigned(35 downto 0);
signal n21 : unsigned(35 downto 0);
signal n22 : unsigned(35 downto 0);
signal n23 : unsigned(35 downto 0);
signal n24 : unsigned(35 downto 0);
signal s25_1 : unsigned(0 downto 0);
signal s26_1 : unsigned(35 downto 0);
signal s26_2 : unsigned(35 downto 0);
signal s27_1 : unsigned(6 downto 0);
signal s27_2 : unsigned(0 downto 0);
signal s28_1 : unsigned(0 downto 0);
signal s28_2 : unsigned(0 downto 0);
signal s28_3 : unsigned(71 downto 0);
signal s29_1 : unsigned(71 downto 0);
component cf_fft_256_18_30 is
port (
clock_c : in std_logic;
i1 : in  unsigned(1 downto 0);
i2 : in  unsigned(0 downto 0);
i3 : in  unsigned(0 downto 0);
o1 : out unsigned(0 downto 0));
end component cf_fft_256_18_30;
component cf_fft_256_18_9 is
port (
clock_c : in std_logic;
i1 : in  unsigned(35 downto 0);
i2 : in  unsigned(35 downto 0);
i3 : in  unsigned(2 downto 0);
i4 : in  unsigned(0 downto 0);
i5 : in  unsigned(0 downto 0);
o1 : out unsigned(35 downto 0);
o2 : out unsigned(35 downto 0));
end component cf_fft_256_18_9;
component cf_fft_256_18_21 is
port (
clock_c : in std_logic;
i1 : in  unsigned(0 downto 0);
i2 : in  unsigned(0 downto 0);
i3 : in  unsigned(0 downto 0);
o1 : out unsigned(6 downto 0);
o2 : out unsigned(0 downto 0));
end component cf_fft_256_18_21;
component cf_fft_256_18_18 is
port (
clock_c : in std_logic;
i1 : in  unsigned(71 downto 0);
i2 : in  unsigned(0 downto 0);
i3 : in  unsigned(5 downto 0);
i4 : in  unsigned(0 downto 0);
i5 : in  unsigned(0 downto 0);
i6 : in  unsigned(0 downto 0);
o1 : out unsigned(0 downto 0);
o2 : out unsigned(0 downto 0);
o3 : out unsigned(71 downto 0));
end component cf_fft_256_18_18;
component cf_fft_256_18_17 is
port (
clock_c : in std_logic;
i1 : in  unsigned(71 downto 0);
i2 : in  unsigned(0 downto 0);
i3 : in  unsigned(5 downto 0);
i4 : in  unsigned(0 downto 0);
i5 : in  unsigned(0 downto 0);
i6 : in  unsigned(0 downto 0);
o1 : out unsigned(71 downto 0));
end component cf_fft_256_18_17;
begin
n1 <= s27_1(6 downto 6) &
  s27_1(5 downto 5) &
  s27_1(4 downto 4);
n2 <= s26_1 & s26_2;
process (clock_c) begin
  if rising_edge(clock_c) then
    if i5 = "1" then
      n3 <= "0";
    elsif i4 = "1" then
      n3 <= s27_2;
    end if;
  end if;
end process;
process (clock_c) begin
  if rising_edge(clock_c) then
    if i5 = "1" then
      n4 <= "0";
    elsif i4 = "1" then
      n4 <= n3;
    end if;
  end if;
end process;
process (clock_c) begin
  if rising_edge(clock_c) then
    if i5 = "1" then
      n5 <= "0";
    elsif i4 = "1" then
      n5 <= n4;
    end if;
  end if;
end process;
process (clock_c) begin
  if rising_edge(clock_c) then
    if i5 = "1" then
      n6 <= "0";
    elsif i4 = "1" then
      n6 <= n5;
    end if;
  end if;
end process;
n7 <= s27_1(6 downto 6) &
  s27_1(5 downto 5) &
  s27_1(4 downto 4) &
  s27_1(3 downto 3) &
  s27_1(2 downto 2) &
  s27_1(1 downto 1);
process (clock_c) begin
  if rising_edge(clock_c) then
    if i5 = "1" then
      n8 <= "000000";
    elsif i4 = "1" then
      n8 <= n7;
    end if;
  end if;
end process;
process (clock_c) begin
  if rising_edge(clock_c) then
    if i5 = "1" then
      n9 <= "000000";
    elsif i4 = "1" then
      n9 <= n8;
    end if;
  end if;
end process;
process (clock_c) begin
  if rising_edge(clock_c) then
    if i5 = "1" then
      n10 <= "000000";
    elsif i4 = "1" then
      n10 <= n9;
    end if;
  end if;
end process;
process (clock_c) begin
  if rising_edge(clock_c) then
    if i5 = "1" then
      n11 <= "000000";
    elsif i4 = "1" then
      n11 <= n10;
    end if;
  end if;
end process;
n12 <= s27_1(0 downto 0);
process (clock_c) begin
  if rising_edge(clock_c) then
    if i5 = "1" then
      n13 <= "0";
    elsif i4 = "1" then
      n13 <= n12;
    end if;
  end if;
end process;
process (clock_c) begin
  if rising_edge(clock_c) then
    if i5 = "1" then
      n14 <= "0";
    elsif i4 = "1" then
      n14 <= n13;
    end if;
  end if;
end process;
process (clock_c) begin
  if rising_edge(clock_c) then
    if i5 = "1" then
      n15 <= "0";
    elsif i4 = "1" then
      n15 <= n14;
    end if;
  end if;
end process;
process (clock_c) begin
  if rising_edge(clock_c) then
    if i5 = "1" then
      n16 <= "0";
    elsif i4 = "1" then
      n16 <= n15;
    end if;
  end if;
end process;
n17 <= not n16;
n18 <= s28_2 & s28_1;
n19 <= s28_3(71 downto 71) &
  s28_3(70 downto 70) &
  s28_3(69 downto 69) &
  s28_3(68 downto 68) &
  s28_3(67 downto 67) &
  s28_3(66 downto 66) &
  s28_3(65 downto 65) &
  s28_3(64 downto 64) &
  s28_3(63 downto 63) &
  s28_3(62 downto 62) &
  s28_3(61 downto 61) &
  s28_3(60 downto 60) &
  s28_3(59 downto 59) &
  s28_3(58 downto 58) &
  s28_3(57 downto 57) &
  s28_3(56 downto 56) &
  s28_3(55 downto 55) &
  s28_3(54 downto 54) &
  s28_3(53 downto 53) &
  s28_3(52 downto 52) &
  s28_3(51 downto 51) &
  s28_3(50 downto 50) &
  s28_3(49 downto 49) &
  s28_3(48 downto 48) &
  s28_3(47 downto 47) &
  s28_3(46 downto 46) &
  s28_3(45 downto 45) &
  s28_3(44 downto 44) &
  s28_3(43 downto 43) &
  s28_3(42 downto 42) &
  s28_3(41 downto 41) &
  s28_3(40 downto 40) &
  s28_3(39 downto 39) &
  s28_3(38 downto 38) &
  s28_3(37 downto 37) &
  s28_3(36 downto 36);
n20 <= s28_3(35 downto 35) &
  s28_3(34 downto 34) &
  s28_3(33 downto 33) &
  s28_3(32 downto 32) &
  s28_3(31 downto 31) &
  s28_3(30 downto 30) &
  s28_3(29 downto 29) &
  s28_3(28 downto 28) &
  s28_3(27 downto 27) &
  s28_3(26 downto 26) &
  s28_3(25 downto 25) &
  s28_3(24 downto 24) &
  s28_3(23 downto 23) &
  s28_3(22 downto 22) &
  s28_3(21 downto 21) &
  s28_3(20 downto 20) &
  s28_3(19 downto 19) &
  s28_3(18 downto 18) &
  s28_3(17 downto 17) &
  s28_3(16 downto 16) &
  s28_3(15 downto 15) &
  s28_3(14 downto 14) &
  s28_3(13 downto 13) &
  s28_3(12 downto 12) &
  s28_3(11 downto 11) &
  s28_3(10 downto 10) &
  s28_3(9 downto 9) &
  s28_3(8 downto 8) &
  s28_3(7 downto 7) &
  s28_3(6 downto 6) &
  s28_3(5 downto 5) &
  s28_3(4 downto 4) &
  s28_3(3 downto 3) &
  s28_3(2 downto 2) &
  s28_3(1 downto 1) &
  s28_3(0 downto 0);
n21 <= s29_1(71 downto 71) &
  s29_1(70 downto 70) &
  s29_1(69 downto 69) &
  s29_1(68 downto 68) &
  s29_1(67 downto 67) &
  s29_1(66 downto 66) &
  s29_1(65 downto 65) &
  s29_1(64 downto 64) &
  s29_1(63 downto 63) &
  s29_1(62 downto 62) &
  s29_1(61 downto 61) &
  s29_1(60 downto 60) &
  s29_1(59 downto 59) &
  s29_1(58 downto 58) &
  s29_1(57 downto 57) &
  s29_1(56 downto 56) &
  s29_1(55 downto 55) &
  s29_1(54 downto 54) &
  s29_1(53 downto 53) &
  s29_1(52 downto 52) &
  s29_1(51 downto 51) &
  s29_1(50 downto 50) &
  s29_1(49 downto 49) &
  s29_1(48 downto 48) &
  s29_1(47 downto 47) &
  s29_1(46 downto 46) &
  s29_1(45 downto 45) &
  s29_1(44 downto 44) &
  s29_1(43 downto 43) &
  s29_1(42 downto 42) &
  s29_1(41 downto 41) &
  s29_1(40 downto 40) &
  s29_1(39 downto 39) &
  s29_1(38 downto 38) &
  s29_1(37 downto 37) &
  s29_1(36 downto 36);
n22 <= s29_1(35 downto 35) &
  s29_1(34 downto 34) &
  s29_1(33 downto 33) &
  s29_1(32 downto 32) &
  s29_1(31 downto 31) &
  s29_1(30 downto 30) &
  s29_1(29 downto 29) &
  s29_1(28 downto 28) &
  s29_1(27 downto 27) &
  s29_1(26 downto 26) &
  s29_1(25 downto 25) &
  s29_1(24 downto 24) &
  s29_1(23 downto 23) &
  s29_1(22 downto 22) &
  s29_1(21 downto 21) &
  s29_1(20 downto 20) &
  s29_1(19 downto 19) &
  s29_1(18 downto 18) &
  s29_1(17 downto 17) &
  s29_1(16 downto 16) &
  s29_1(15 downto 15) &
  s29_1(14 downto 14) &
  s29_1(13 downto 13) &
  s29_1(12 downto 12) &
  s29_1(11 downto 11) &
  s29_1(10 downto 10) &
  s29_1(9 downto 9) &
  s29_1(8 downto 8) &
  s29_1(7 downto 7) &
  s29_1(6 downto 6) &
  s29_1(5 downto 5) &
  s29_1(4 downto 4) &
  s29_1(3 downto 3) &
  s29_1(2 downto 2) &
  s29_1(1 downto 1) &
  s29_1(0 downto 0);
n23 <= n20 when s25_1 = "1" else n19;
n24 <= n22 when s25_1 = "1" else n21;
s25 : cf_fft_256_18_30 port map (clock_c, n18, i4, i5, s25_1);
s26 : cf_fft_256_18_9 port map (clock_c, i2, i3, n1, i4, i5, s26_1, s26_2);
s27 : cf_fft_256_18_21 port map (clock_c, i1, i4, i5, s27_1, s27_2);
s28 : cf_fft_256_18_18 port map (clock_c, n2, n6, n11, n17, i4, i5, s28_1, s28_2, s28_3);
s29 : cf_fft_256_18_17 port map (clock_c, n2, n6, n11, n16, i4, i5, s29_1);
o3 <= n24;
o2 <= n23;
o1 <= s28_1;
end architecture rtl;

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
entity cf_fft_256_18_7 is
port (
clock_c : in std_logic;
i1 : in  unsigned(35 downto 0);
i2 : in  unsigned(35 downto 0);
i3 : in  unsigned(1 downto 0);
i4 : in  unsigned(0 downto 0);
i5 : in  unsigned(0 downto 0);
o1 : out unsigned(35 downto 0);
o2 : out unsigned(35 downto 0));
end entity cf_fft_256_18_7;
architecture rtl of cf_fft_256_18_7 is
signal n1 : unsigned(35 downto 0) := "000000000000000000000000000000000000";
signal n2 : unsigned(17 downto 0);
signal n3 : unsigned(17 downto 0);
signal n4 : unsigned(35 downto 0) := "000000000000000000000000000000000000";
signal n5 : unsigned(17 downto 0);
signal n6 : unsigned(17 downto 0);
signal n7 : unsigned(17 downto 0) := "000000000000000000";
signal n8 : unsigned(17 downto 0) := "000000000000000000";
signal n9 : unsigned(17 downto 0) := "000000000000000000";
signal n10 : unsigned(17 downto 0) := "000000000000000000";
signal n11 : unsigned(35 downto 0) := "000000000000000000000000000000000000";
signal n12 : unsigned(17 downto 0);
signal n13 : unsigned(17 downto 0);
signal n14 : unsigned(35 downto 0);
signal n15 : unsigned(17 downto 0);
signal n16 : unsigned(17 downto 0) := "000000000000000000";
signal n17 : unsigned(35 downto 0);
signal n18 : unsigned(17 downto 0);
signal n19 : unsigned(17 downto 0) := "000000000000000000";
signal n20 : unsigned(17 downto 0);
signal n21 : unsigned(17 downto 0) := "000000000000000000";
signal n22 : unsigned(35 downto 0);
signal n23 : unsigned(17 downto 0);
signal n24 : unsigned(17 downto 0) := "000000000000000000";
signal n25 : unsigned(35 downto 0);
signal n26 : unsigned(17 downto 0);
signal n27 : unsigned(17 downto 0) := "000000000000000000";
signal n28 : unsigned(17 downto 0);
signal n29 : unsigned(17 downto 0) := "000000000000000000";
signal n30 : unsigned(17 downto 0);
signal n31 : unsigned(17 downto 0);
signal n32 : unsigned(35 downto 0);
signal n33 : unsigned(35 downto 0) := "000000000000000000000000000000000000";
signal n34 : unsigned(17 downto 0);
signal n35 : unsigned(17 downto 0);
signal n36 : unsigned(35 downto 0);
signal n37 : unsigned(35 downto 0) := "000000000000000000000000000000000000";
begin
process (clock_c) begin
  if rising_edge(clock_c) then
    if i5 = "1" then
      n1 <= "000000000000000000000000000000000000";
    elsif i4 = "1" then
      n1 <= i1;
    end if;
  end if;
end process;
n2 <= n1(35 downto 35) &
  n1(34 downto 34) &
  n1(33 downto 33) &
  n1(32 downto 32) &
  n1(31 downto 31) &
  n1(30 downto 30) &
  n1(29 downto 29) &
  n1(28 downto 28) &
  n1(27 downto 27) &
  n1(26 downto 26) &
  n1(25 downto 25) &
  n1(24 downto 24) &
  n1(23 downto 23) &
  n1(22 downto 22) &
  n1(21 downto 21) &
  n1(20 downto 20) &
  n1(19 downto 19) &
  n1(18 downto 18);
n3 <= n1(17 downto 17) &
  n1(16 downto 16) &
  n1(15 downto 15) &
  n1(14 downto 14) &
  n1(13 downto 13) &
  n1(12 downto 12) &
  n1(11 downto 11) &
  n1(10 downto 10) &
  n1(9 downto 9) &
  n1(8 downto 8) &
  n1(7 downto 7) &
  n1(6 downto 6) &
  n1(5 downto 5) &
  n1(4 downto 4) &
  n1(3 downto 3) &
  n1(2 downto 2) &
  n1(1 downto 1) &
  n1(0 downto 0);
process (clock_c) begin
  if rising_edge(clock_c) then
    if i5 = "1" then
      n4 <= "000000000000000000000000000000000000";
    elsif i4 = "1" then
      n4 <= i2;
    end if;
  end if;
end process;
n5 <= n4(35 downto 35) &
  n4(34 downto 34) &
  n4(33 downto 33) &
  n4(32 downto 32) &
  n4(31 downto 31) &
  n4(30 downto 30) &
  n4(29 downto 29) &
  n4(28 downto 28) &
  n4(27 downto 27) &
  n4(26 downto 26) &
  n4(25 downto 25) &
  n4(24 downto 24) &
  n4(23 downto 23) &
  n4(22 downto 22) &
  n4(21 downto 21) &
  n4(20 downto 20) &
  n4(19 downto 19) &
  n4(18 downto 18);
n6 <= n4(17 downto 17) &
  n4(16 downto 16) &
  n4(15 downto 15) &
  n4(14 downto 14) &
  n4(13 downto 13) &
  n4(12 downto 12) &
  n4(11 downto 11) &
  n4(10 downto 10) &
  n4(9 downto 9) &
  n4(8 downto 8) &
  n4(7 downto 7) &
  n4(6 downto 6) &
  n4(5 downto 5) &
  n4(4 downto 4) &
  n4(3 downto 3) &
  n4(2 downto 2) &
  n4(1 downto 1) &
  n4(0 downto 0);
process (clock_c) begin
  if rising_edge(clock_c) then
    if i5 = "1" then
      n7 <= "000000000000000000";
    elsif i4 = "1" then
      n7 <= n2;
    end if;
  end if;
end process;
process (clock_c) begin
  if rising_edge(clock_c) then
    if i5 = "1" then
      n8 <= "000000000000000000";
    elsif i4 = "1" then
      n8 <= n7;
    end if;
  end if;
end process;
process (clock_c) begin
  if rising_edge(clock_c) then
    if i5 = "1" then
      n9 <= "000000000000000000";
    elsif i4 = "1" then
      n9 <= n3;
    end if;
  end if;
end process;
process (clock_c) begin
  if rising_edge(clock_c) then
    if i5 = "1" then
      n10 <= "000000000000000000";
    elsif i4 = "1" then
      n10 <= n9;
    end if;
  end if;
end process;
process (clock_c) begin
  if rising_edge(clock_c) then 
    if i4 = "1" then
      case i3 is
        when "00" => n11 <= "011111111111111111000000000000000000";
        when "01" => n11 <= "010110101000001001101001010111110110";
        when "10" => n11 <= "000000000000000000100000000000000000";
        when "11" => n11 <= "101001010111110110101001010111110110";
        when others => n11 <= "XXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX";
      end case;
    end if;
  end if;
end process;
n12 <= n11(35 downto 35) &
  n11(34 downto 34) &
  n11(33 downto 33) &
  n11(32 downto 32) &
  n11(31 downto 31) &
  n11(30 downto 30) &
  n11(29 downto 29) &
  n11(28 downto 28) &
  n11(27 downto 27) &
  n11(26 downto 26) &
  n11(25 downto 25) &
  n11(24 downto 24) &
  n11(23 downto 23) &
  n11(22 downto 22) &
  n11(21 downto 21) &
  n11(20 downto 20) &
  n11(19 downto 19) &
  n11(18 downto 18);
n13 <= n11(17 downto 17) &
  n11(16 downto 16) &
  n11(15 downto 15) &
  n11(14 downto 14) &
  n11(13 downto 13) &
  n11(12 downto 12) &
  n11(11 downto 11) &
  n11(10 downto 10) &
  n11(9 downto 9) &
  n11(8 downto 8) &
  n11(7 downto 7) &
  n11(6 downto 6) &
  n11(5 downto 5) &
  n11(4 downto 4) &
  n11(3 downto 3) &
  n11(2 downto 2) &
  n11(1 downto 1) &
  n11(0 downto 0);
n14 <= unsigned(signed(n5) * signed(n12));
n15 <= n14(34 downto 34) &
  n14(33 downto 33) &
  n14(32 downto 32) &
  n14(31 downto 31) &
  n14(30 downto 30) &
  n14(29 downto 29) &
  n14(28 downto 28) &
  n14(27 downto 27) &
  n14(26 downto 26) &
  n14(25 downto 25) &
  n14(24 downto 24) &
  n14(23 downto 23) &
  n14(22 downto 22) &
  n14(21 downto 21) &
  n14(20 downto 20) &
  n14(19 downto 19) &
  n14(18 downto 18) &
  n14(17 downto 17);
process (clock_c) begin
  if rising_edge(clock_c) then
    if i5 = "1" then
      n16 <= "000000000000000000";
    elsif i4 = "1" then
      n16 <= n15;
    end if;
  end if;
end process;
n17 <= unsigned(signed(n6) * signed(n13));
n18 <= n17(34 downto 34) &
  n17(33 downto 33) &
  n17(32 downto 32) &
  n17(31 downto 31) &
  n17(30 downto 30) &
  n17(29 downto 29) &
  n17(28 downto 28) &
  n17(27 downto 27) &
  n17(26 downto 26) &
  n17(25 downto 25) &
  n17(24 downto 24) &
  n17(23 downto 23) &
  n17(22 downto 22) &
  n17(21 downto 21) &
  n17(20 downto 20) &
  n17(19 downto 19) &
  n17(18 downto 18) &
  n17(17 downto 17);
process (clock_c) begin
  if rising_edge(clock_c) then
    if i5 = "1" then
      n19 <= "000000000000000000";
    elsif i4 = "1" then
      n19 <= n18;
    end if;
  end if;
end process;
n20 <= n16 - n19;
process (clock_c) begin
  if rising_edge(clock_c) then
    if i5 = "1" then
      n21 <= "000000000000000000";
    elsif i4 = "1" then
      n21 <= n20;
    end if;
  end if;
end process;
n22 <= unsigned(signed(n5) * signed(n13));
n23 <= n22(34 downto 34) &
  n22(33 downto 33) &
  n22(32 downto 32) &
  n22(31 downto 31) &
  n22(30 downto 30) &
  n22(29 downto 29) &
  n22(28 downto 28) &
  n22(27 downto 27) &
  n22(26 downto 26) &
  n22(25 downto 25) &
  n22(24 downto 24) &
  n22(23 downto 23) &
  n22(22 downto 22) &
  n22(21 downto 21) &
  n22(20 downto 20) &
  n22(19 downto 19) &
  n22(18 downto 18) &
  n22(17 downto 17);
process (clock_c) begin
  if rising_edge(clock_c) then
    if i5 = "1" then
      n24 <= "000000000000000000";
    elsif i4 = "1" then
      n24 <= n23;
    end if;
  end if;
end process;
n25 <= unsigned(signed(n6) * signed(n12));
n26 <= n25(34 downto 34) &
  n25(33 downto 33) &
  n25(32 downto 32) &
  n25(31 downto 31) &
  n25(30 downto 30) &
  n25(29 downto 29) &
  n25(28 downto 28) &
  n25(27 downto 27) &
  n25(26 downto 26) &
  n25(25 downto 25) &
  n25(24 downto 24) &
  n25(23 downto 23) &
  n25(22 downto 22) &
  n25(21 downto 21) &
  n25(20 downto 20) &
  n25(19 downto 19) &
  n25(18 downto 18) &
  n25(17 downto 17);
process (clock_c) begin
  if rising_edge(clock_c) then
    if i5 = "1" then
      n27 <= "000000000000000000";
    elsif i4 = "1" then
      n27 <= n26;
    end if;
  end if;
end process;
n28 <= n24 + n27;
process (clock_c) begin
  if rising_edge(clock_c) then
    if i5 = "1" then
      n29 <= "000000000000000000";
    elsif i4 = "1" then
      n29 <= n28;
    end if;
  end if;
end process;
n30 <= n8 + n21;
n31 <= n10 + n29;
n32 <= n30 & n31;
process (clock_c) begin
  if rising_edge(clock_c) then
    if i5 = "1" then
      n33 <= "000000000000000000000000000000000000";
    elsif i4 = "1" then
      n33 <= n32;
    end if;
  end if;
end process;
n34 <= n8 - n21;
n35 <= n10 - n29;
n36 <= n34 & n35;
process (clock_c) begin
  if rising_edge(clock_c) then
    if i5 = "1" then
      n37 <= "000000000000000000000000000000000000";
    elsif i4 = "1" then
      n37 <= n36;
    end if;
  end if;
end process;
o2 <= n37;
o1 <= n33;
end architecture rtl;

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
entity cf_fft_256_18_6 is
port (
clock_c : in std_logic;
i1 : in  unsigned(0 downto 0);
i2 : in  unsigned(35 downto 0);
i3 : in  unsigned(35 downto 0);
i4 : in  unsigned(0 downto 0);
i5 : in  unsigned(0 downto 0);
o1 : out unsigned(0 downto 0);
o2 : out unsigned(35 downto 0);
o3 : out unsigned(35 downto 0));
end entity cf_fft_256_18_6;
architecture rtl of cf_fft_256_18_6 is
signal n1 : unsigned(1 downto 0);
signal n2 : unsigned(71 downto 0);
signal n3 : unsigned(0 downto 0) := "0";
signal n4 : unsigned(0 downto 0) := "0";
signal n5 : unsigned(0 downto 0) := "0";
signal n6 : unsigned(0 downto 0) := "0";
signal n7 : unsigned(5 downto 0);
signal n8 : unsigned(5 downto 0) := "000000";
signal n9 : unsigned(5 downto 0) := "000000";
signal n10 : unsigned(5 downto 0) := "000000";
signal n11 : unsigned(5 downto 0) := "000000";
signal n12 : unsigned(0 downto 0);
signal n13 : unsigned(0 downto 0) := "0";
signal n14 : unsigned(0 downto 0) := "0";
signal n15 : unsigned(0 downto 0) := "0";
signal n16 : unsigned(0 downto 0) := "0";
signal n17 : unsigned(0 downto 0);
signal n18 : unsigned(1 downto 0);
signal n19 : unsigned(35 downto 0);
signal n20 : unsigned(35 downto 0);
signal n21 : unsigned(35 downto 0);
signal n22 : unsigned(35 downto 0);
signal n23 : unsigned(35 downto 0);
signal n24 : unsigned(35 downto 0);
signal s25_1 : unsigned(0 downto 0);
signal s26_1 : unsigned(35 downto 0);
signal s26_2 : unsigned(35 downto 0);
signal s27_1 : unsigned(6 downto 0);
signal s27_2 : unsigned(0 downto 0);
signal s28_1 : unsigned(0 downto 0);
signal s28_2 : unsigned(0 downto 0);
signal s28_3 : unsigned(71 downto 0);
signal s29_1 : unsigned(71 downto 0);
component cf_fft_256_18_30 is
port (
clock_c : in std_logic;
i1 : in  unsigned(1 downto 0);
i2 : in  unsigned(0 downto 0);
i3 : in  unsigned(0 downto 0);
o1 : out unsigned(0 downto 0));
end component cf_fft_256_18_30;
component cf_fft_256_18_7 is
port (
clock_c : in std_logic;
i1 : in  unsigned(35 downto 0);
i2 : in  unsigned(35 downto 0);
i3 : in  unsigned(1 downto 0);
i4 : in  unsigned(0 downto 0);
i5 : in  unsigned(0 downto 0);
o1 : out unsigned(35 downto 0);
o2 : out unsigned(35 downto 0));
end component cf_fft_256_18_7;
component cf_fft_256_18_21 is
port (
clock_c : in std_logic;
i1 : in  unsigned(0 downto 0);
i2 : in  unsigned(0 downto 0);
i3 : in  unsigned(0 downto 0);
o1 : out unsigned(6 downto 0);
o2 : out unsigned(0 downto 0));
end component cf_fft_256_18_21;
component cf_fft_256_18_18 is
port (
clock_c : in std_logic;
i1 : in  unsigned(71 downto 0);
i2 : in  unsigned(0 downto 0);
i3 : in  unsigned(5 downto 0);
i4 : in  unsigned(0 downto 0);
i5 : in  unsigned(0 downto 0);
i6 : in  unsigned(0 downto 0);
o1 : out unsigned(0 downto 0);
o2 : out unsigned(0 downto 0);
o3 : out unsigned(71 downto 0));
end component cf_fft_256_18_18;
component cf_fft_256_18_17 is
port (
clock_c : in std_logic;
i1 : in  unsigned(71 downto 0);
i2 : in  unsigned(0 downto 0);
i3 : in  unsigned(5 downto 0);
i4 : in  unsigned(0 downto 0);
i5 : in  unsigned(0 downto 0);
i6 : in  unsigned(0 downto 0);
o1 : out unsigned(71 downto 0));
end component cf_fft_256_18_17;
begin
n1 <= s27_1(6 downto 6) &
  s27_1(5 downto 5);
n2 <= s26_1 & s26_2;
process (clock_c) begin
  if rising_edge(clock_c) then
    if i5 = "1" then
      n3 <= "0";
    elsif i4 = "1" then
      n3 <= s27_2;
    end if;
  end if;
end process;
process (clock_c) begin
  if rising_edge(clock_c) then
    if i5 = "1" then
      n4 <= "0";
    elsif i4 = "1" then
      n4 <= n3;
    end if;
  end if;
end process;
process (clock_c) begin
  if rising_edge(clock_c) then
    if i5 = "1" then
      n5 <= "0";
    elsif i4 = "1" then
      n5 <= n4;
    end if;
  end if;
end process;
process (clock_c) begin
  if rising_edge(clock_c) then
    if i5 = "1" then
      n6 <= "0";
    elsif i4 = "1" then
      n6 <= n5;
    end if;
  end if;
end process;
n7 <= s27_1(6 downto 6) &
  s27_1(5 downto 5) &
  s27_1(4 downto 4) &
  s27_1(3 downto 3) &
  s27_1(2 downto 2) &
  s27_1(1 downto 1);
process (clock_c) begin
  if rising_edge(clock_c) then
    if i5 = "1" then
      n8 <= "000000";
    elsif i4 = "1" then
      n8 <= n7;
    end if;
  end if;
end process;
process (clock_c) begin
  if rising_edge(clock_c) then
    if i5 = "1" then
      n9 <= "000000";
    elsif i4 = "1" then
      n9 <= n8;
    end if;
  end if;
end process;
process (clock_c) begin
  if rising_edge(clock_c) then
    if i5 = "1" then
      n10 <= "000000";
    elsif i4 = "1" then
      n10 <= n9;
    end if;
  end if;
end process;
process (clock_c) begin
  if rising_edge(clock_c) then
    if i5 = "1" then
      n11 <= "000000";
    elsif i4 = "1" then
      n11 <= n10;
    end if;
  end if;
end process;
n12 <= s27_1(0 downto 0);
process (clock_c) begin
  if rising_edge(clock_c) then
    if i5 = "1" then
      n13 <= "0";
    elsif i4 = "1" then
      n13 <= n12;
    end if;
  end if;
end process;
process (clock_c) begin
  if rising_edge(clock_c) then
    if i5 = "1" then
      n14 <= "0";
    elsif i4 = "1" then
      n14 <= n13;
    end if;
  end if;
end process;
process (clock_c) begin
  if rising_edge(clock_c) then
    if i5 = "1" then
      n15 <= "0";
    elsif i4 = "1" then
      n15 <= n14;
    end if;
  end if;
end process;
process (clock_c) begin
  if rising_edge(clock_c) then
    if i5 = "1" then
      n16 <= "0";
    elsif i4 = "1" then
      n16 <= n15;
    end if;
  end if;
end process;
n17 <= not n16;
n18 <= s28_2 & s28_1;
n19 <= s28_3(71 downto 71) &
  s28_3(70 downto 70) &
  s28_3(69 downto 69) &
  s28_3(68 downto 68) &
  s28_3(67 downto 67) &
  s28_3(66 downto 66) &
  s28_3(65 downto 65) &
  s28_3(64 downto 64) &
  s28_3(63 downto 63) &
  s28_3(62 downto 62) &
  s28_3(61 downto 61) &
  s28_3(60 downto 60) &
  s28_3(59 downto 59) &
  s28_3(58 downto 58) &
  s28_3(57 downto 57) &
  s28_3(56 downto 56) &
  s28_3(55 downto 55) &
  s28_3(54 downto 54) &
  s28_3(53 downto 53) &
  s28_3(52 downto 52) &
  s28_3(51 downto 51) &
  s28_3(50 downto 50) &
  s28_3(49 downto 49) &
  s28_3(48 downto 48) &
  s28_3(47 downto 47) &
  s28_3(46 downto 46) &
  s28_3(45 downto 45) &
  s28_3(44 downto 44) &
  s28_3(43 downto 43) &
  s28_3(42 downto 42) &
  s28_3(41 downto 41) &
  s28_3(40 downto 40) &
  s28_3(39 downto 39) &
  s28_3(38 downto 38) &
  s28_3(37 downto 37) &
  s28_3(36 downto 36);
n20 <= s28_3(35 downto 35) &
  s28_3(34 downto 34) &
  s28_3(33 downto 33) &
  s28_3(32 downto 32) &
  s28_3(31 downto 31) &
  s28_3(30 downto 30) &
  s28_3(29 downto 29) &
  s28_3(28 downto 28) &
  s28_3(27 downto 27) &
  s28_3(26 downto 26) &
  s28_3(25 downto 25) &
  s28_3(24 downto 24) &
  s28_3(23 downto 23) &
  s28_3(22 downto 22) &
  s28_3(21 downto 21) &
  s28_3(20 downto 20) &
  s28_3(19 downto 19) &
  s28_3(18 downto 18) &
  s28_3(17 downto 17) &
  s28_3(16 downto 16) &
  s28_3(15 downto 15) &
  s28_3(14 downto 14) &
  s28_3(13 downto 13) &
  s28_3(12 downto 12) &
  s28_3(11 downto 11) &
  s28_3(10 downto 10) &
  s28_3(9 downto 9) &
  s28_3(8 downto 8) &
  s28_3(7 downto 7) &
  s28_3(6 downto 6) &
  s28_3(5 downto 5) &
  s28_3(4 downto 4) &
  s28_3(3 downto 3) &
  s28_3(2 downto 2) &
  s28_3(1 downto 1) &
  s28_3(0 downto 0);
n21 <= s29_1(71 downto 71) &
  s29_1(70 downto 70) &
  s29_1(69 downto 69) &
  s29_1(68 downto 68) &
  s29_1(67 downto 67) &
  s29_1(66 downto 66) &
  s29_1(65 downto 65) &
  s29_1(64 downto 64) &
  s29_1(63 downto 63) &
  s29_1(62 downto 62) &
  s29_1(61 downto 61) &
  s29_1(60 downto 60) &
  s29_1(59 downto 59) &
  s29_1(58 downto 58) &
  s29_1(57 downto 57) &
  s29_1(56 downto 56) &
  s29_1(55 downto 55) &
  s29_1(54 downto 54) &
  s29_1(53 downto 53) &
  s29_1(52 downto 52) &
  s29_1(51 downto 51) &
  s29_1(50 downto 50) &
  s29_1(49 downto 49) &
  s29_1(48 downto 48) &
  s29_1(47 downto 47) &
  s29_1(46 downto 46) &
  s29_1(45 downto 45) &
  s29_1(44 downto 44) &
  s29_1(43 downto 43) &
  s29_1(42 downto 42) &
  s29_1(41 downto 41) &
  s29_1(40 downto 40) &
  s29_1(39 downto 39) &
  s29_1(38 downto 38) &
  s29_1(37 downto 37) &
  s29_1(36 downto 36);
n22 <= s29_1(35 downto 35) &
  s29_1(34 downto 34) &
  s29_1(33 downto 33) &
  s29_1(32 downto 32) &
  s29_1(31 downto 31) &
  s29_1(30 downto 30) &
  s29_1(29 downto 29) &
  s29_1(28 downto 28) &
  s29_1(27 downto 27) &
  s29_1(26 downto 26) &
  s29_1(25 downto 25) &
  s29_1(24 downto 24) &
  s29_1(23 downto 23) &
  s29_1(22 downto 22) &
  s29_1(21 downto 21) &
  s29_1(20 downto 20) &
  s29_1(19 downto 19) &
  s29_1(18 downto 18) &
  s29_1(17 downto 17) &
  s29_1(16 downto 16) &
  s29_1(15 downto 15) &
  s29_1(14 downto 14) &
  s29_1(13 downto 13) &
  s29_1(12 downto 12) &
  s29_1(11 downto 11) &
  s29_1(10 downto 10) &
  s29_1(9 downto 9) &
  s29_1(8 downto 8) &
  s29_1(7 downto 7) &
  s29_1(6 downto 6) &
  s29_1(5 downto 5) &
  s29_1(4 downto 4) &
  s29_1(3 downto 3) &
  s29_1(2 downto 2) &
  s29_1(1 downto 1) &
  s29_1(0 downto 0);
n23 <= n20 when s25_1 = "1" else n19;
n24 <= n22 when s25_1 = "1" else n21;
s25 : cf_fft_256_18_30 port map (clock_c, n18, i4, i5, s25_1);
s26 : cf_fft_256_18_7 port map (clock_c, i2, i3, n1, i4, i5, s26_1, s26_2);
s27 : cf_fft_256_18_21 port map (clock_c, i1, i4, i5, s27_1, s27_2);
s28 : cf_fft_256_18_18 port map (clock_c, n2, n6, n11, n17, i4, i5, s28_1, s28_2, s28_3);
s29 : cf_fft_256_18_17 port map (clock_c, n2, n6, n11, n16, i4, i5, s29_1);
o3 <= n24;
o2 <= n23;
o1 <= s28_1;
end architecture rtl;

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
entity cf_fft_256_18_5 is
port (
clock_c : in std_logic;
i1 : in  unsigned(35 downto 0);
i2 : in  unsigned(35 downto 0);
i3 : in  unsigned(0 downto 0);
i4 : in  unsigned(0 downto 0);
i5 : in  unsigned(0 downto 0);
o1 : out unsigned(35 downto 0);
o2 : out unsigned(35 downto 0));
end entity cf_fft_256_18_5;
architecture rtl of cf_fft_256_18_5 is
signal n1 : unsigned(35 downto 0) := "000000000000000000000000000000000000";
signal n2 : unsigned(17 downto 0);
signal n3 : unsigned(17 downto 0);
signal n4 : unsigned(35 downto 0) := "000000000000000000000000000000000000";
signal n5 : unsigned(17 downto 0);
signal n6 : unsigned(17 downto 0);
signal n7 : unsigned(17 downto 0) := "000000000000000000";
signal n8 : unsigned(17 downto 0) := "000000000000000000";
signal n9 : unsigned(17 downto 0) := "000000000000000000";
signal n10 : unsigned(17 downto 0) := "000000000000000000";
signal n11 : unsigned(35 downto 0) := "000000000000000000000000000000000000";
signal n12 : unsigned(17 downto 0);
signal n13 : unsigned(17 downto 0);
signal n14 : unsigned(35 downto 0);
signal n15 : unsigned(17 downto 0);
signal n16 : unsigned(17 downto 0) := "000000000000000000";
signal n17 : unsigned(35 downto 0);
signal n18 : unsigned(17 downto 0);
signal n19 : unsigned(17 downto 0) := "000000000000000000";
signal n20 : unsigned(17 downto 0);
signal n21 : unsigned(17 downto 0) := "000000000000000000";
signal n22 : unsigned(35 downto 0);
signal n23 : unsigned(17 downto 0);
signal n24 : unsigned(17 downto 0) := "000000000000000000";
signal n25 : unsigned(35 downto 0);
signal n26 : unsigned(17 downto 0);
signal n27 : unsigned(17 downto 0) := "000000000000000000";
signal n28 : unsigned(17 downto 0);
signal n29 : unsigned(17 downto 0) := "000000000000000000";
signal n30 : unsigned(17 downto 0);
signal n31 : unsigned(17 downto 0);
signal n32 : unsigned(35 downto 0);
signal n33 : unsigned(35 downto 0) := "000000000000000000000000000000000000";
signal n34 : unsigned(17 downto 0);
signal n35 : unsigned(17 downto 0);
signal n36 : unsigned(35 downto 0);
signal n37 : unsigned(35 downto 0) := "000000000000000000000000000000000000";
begin
process (clock_c) begin
  if rising_edge(clock_c) then
    if i5 = "1" then
      n1 <= "000000000000000000000000000000000000";
    elsif i4 = "1" then
      n1 <= i1;
    end if;
  end if;
end process;
n2 <= n1(35 downto 35) &
  n1(34 downto 34) &
  n1(33 downto 33) &
  n1(32 downto 32) &
  n1(31 downto 31) &
  n1(30 downto 30) &
  n1(29 downto 29) &
  n1(28 downto 28) &
  n1(27 downto 27) &
  n1(26 downto 26) &
  n1(25 downto 25) &
  n1(24 downto 24) &
  n1(23 downto 23) &
  n1(22 downto 22) &
  n1(21 downto 21) &
  n1(20 downto 20) &
  n1(19 downto 19) &
  n1(18 downto 18);
n3 <= n1(17 downto 17) &
  n1(16 downto 16) &
  n1(15 downto 15) &
  n1(14 downto 14) &
  n1(13 downto 13) &
  n1(12 downto 12) &
  n1(11 downto 11) &
  n1(10 downto 10) &
  n1(9 downto 9) &
  n1(8 downto 8) &
  n1(7 downto 7) &
  n1(6 downto 6) &
  n1(5 downto 5) &
  n1(4 downto 4) &
  n1(3 downto 3) &
  n1(2 downto 2) &
  n1(1 downto 1) &
  n1(0 downto 0);
process (clock_c) begin
  if rising_edge(clock_c) then
    if i5 = "1" then
      n4 <= "000000000000000000000000000000000000";
    elsif i4 = "1" then
      n4 <= i2;
    end if;
  end if;
end process;
n5 <= n4(35 downto 35) &
  n4(34 downto 34) &
  n4(33 downto 33) &
  n4(32 downto 32) &
  n4(31 downto 31) &
  n4(30 downto 30) &
  n4(29 downto 29) &
  n4(28 downto 28) &
  n4(27 downto 27) &
  n4(26 downto 26) &
  n4(25 downto 25) &
  n4(24 downto 24) &
  n4(23 downto 23) &
  n4(22 downto 22) &
  n4(21 downto 21) &
  n4(20 downto 20) &
  n4(19 downto 19) &
  n4(18 downto 18);
n6 <= n4(17 downto 17) &
  n4(16 downto 16) &
  n4(15 downto 15) &
  n4(14 downto 14) &
  n4(13 downto 13) &
  n4(12 downto 12) &
  n4(11 downto 11) &
  n4(10 downto 10) &
  n4(9 downto 9) &
  n4(8 downto 8) &
  n4(7 downto 7) &
  n4(6 downto 6) &
  n4(5 downto 5) &
  n4(4 downto 4) &
  n4(3 downto 3) &
  n4(2 downto 2) &
  n4(1 downto 1) &
  n4(0 downto 0);
process (clock_c) begin
  if rising_edge(clock_c) then
    if i5 = "1" then
      n7 <= "000000000000000000";
    elsif i4 = "1" then
      n7 <= n2;
    end if;
  end if;
end process;
process (clock_c) begin
  if rising_edge(clock_c) then
    if i5 = "1" then
      n8 <= "000000000000000000";
    elsif i4 = "1" then
      n8 <= n7;
    end if;
  end if;
end process;
process (clock_c) begin
  if rising_edge(clock_c) then
    if i5 = "1" then
      n9 <= "000000000000000000";
    elsif i4 = "1" then
      n9 <= n3;
    end if;
  end if;
end process;
process (clock_c) begin
  if rising_edge(clock_c) then
    if i5 = "1" then
      n10 <= "000000000000000000";
    elsif i4 = "1" then
      n10 <= n9;
    end if;
  end if;
end process;
process (clock_c) begin
  if rising_edge(clock_c) then 
    if i4 = "1" then
      case i3 is
        when "0" => n11 <= "011111111111111111000000000000000000";
        when "1" => n11 <= "000000000000000000100000000000000000";
        when others => n11 <= "XXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX";
      end case;
    end if;
  end if;
end process;
n12 <= n11(35 downto 35) &
  n11(34 downto 34) &
  n11(33 downto 33) &
  n11(32 downto 32) &
  n11(31 downto 31) &
  n11(30 downto 30) &
  n11(29 downto 29) &
  n11(28 downto 28) &
  n11(27 downto 27) &
  n11(26 downto 26) &
  n11(25 downto 25) &
  n11(24 downto 24) &
  n11(23 downto 23) &
  n11(22 downto 22) &
  n11(21 downto 21) &
  n11(20 downto 20) &
  n11(19 downto 19) &
  n11(18 downto 18);
n13 <= n11(17 downto 17) &
  n11(16 downto 16) &
  n11(15 downto 15) &
  n11(14 downto 14) &
  n11(13 downto 13) &
  n11(12 downto 12) &
  n11(11 downto 11) &
  n11(10 downto 10) &
  n11(9 downto 9) &
  n11(8 downto 8) &
  n11(7 downto 7) &
  n11(6 downto 6) &
  n11(5 downto 5) &
  n11(4 downto 4) &
  n11(3 downto 3) &
  n11(2 downto 2) &
  n11(1 downto 1) &
  n11(0 downto 0);
n14 <= unsigned(signed(n5) * signed(n12));
n15 <= n14(34 downto 34) &
  n14(33 downto 33) &
  n14(32 downto 32) &
  n14(31 downto 31) &
  n14(30 downto 30) &
  n14(29 downto 29) &
  n14(28 downto 28) &
  n14(27 downto 27) &
  n14(26 downto 26) &
  n14(25 downto 25) &
  n14(24 downto 24) &
  n14(23 downto 23) &
  n14(22 downto 22) &
  n14(21 downto 21) &
  n14(20 downto 20) &
  n14(19 downto 19) &
  n14(18 downto 18) &
  n14(17 downto 17);
process (clock_c) begin
  if rising_edge(clock_c) then
    if i5 = "1" then
      n16 <= "000000000000000000";
    elsif i4 = "1" then
      n16 <= n15;
    end if;
  end if;
end process;
n17 <= unsigned(signed(n6) * signed(n13));
n18 <= n17(34 downto 34) &
  n17(33 downto 33) &
  n17(32 downto 32) &
  n17(31 downto 31) &
  n17(30 downto 30) &
  n17(29 downto 29) &
  n17(28 downto 28) &
  n17(27 downto 27) &
  n17(26 downto 26) &
  n17(25 downto 25) &
  n17(24 downto 24) &
  n17(23 downto 23) &
  n17(22 downto 22) &
  n17(21 downto 21) &
  n17(20 downto 20) &
  n17(19 downto 19) &
  n17(18 downto 18) &
  n17(17 downto 17);
process (clock_c) begin
  if rising_edge(clock_c) then
    if i5 = "1" then
      n19 <= "000000000000000000";
    elsif i4 = "1" then
      n19 <= n18;
    end if;
  end if;
end process;
n20 <= n16 - n19;
process (clock_c) begin
  if rising_edge(clock_c) then
    if i5 = "1" then
      n21 <= "000000000000000000";
    elsif i4 = "1" then
      n21 <= n20;
    end if;
  end if;
end process;
n22 <= unsigned(signed(n5) * signed(n13));
n23 <= n22(34 downto 34) &
  n22(33 downto 33) &
  n22(32 downto 32) &
  n22(31 downto 31) &
  n22(30 downto 30) &
  n22(29 downto 29) &
  n22(28 downto 28) &
  n22(27 downto 27) &
  n22(26 downto 26) &
  n22(25 downto 25) &
  n22(24 downto 24) &
  n22(23 downto 23) &
  n22(22 downto 22) &
  n22(21 downto 21) &
  n22(20 downto 20) &
  n22(19 downto 19) &
  n22(18 downto 18) &
  n22(17 downto 17);
process (clock_c) begin
  if rising_edge(clock_c) then
    if i5 = "1" then
      n24 <= "000000000000000000";
    elsif i4 = "1" then
      n24 <= n23;
    end if;
  end if;
end process;
n25 <= unsigned(signed(n6) * signed(n12));
n26 <= n25(34 downto 34) &
  n25(33 downto 33) &
  n25(32 downto 32) &
  n25(31 downto 31) &
  n25(30 downto 30) &
  n25(29 downto 29) &
  n25(28 downto 28) &
  n25(27 downto 27) &
  n25(26 downto 26) &
  n25(25 downto 25) &
  n25(24 downto 24) &
  n25(23 downto 23) &
  n25(22 downto 22) &
  n25(21 downto 21) &
  n25(20 downto 20) &
  n25(19 downto 19) &
  n25(18 downto 18) &
  n25(17 downto 17);
process (clock_c) begin
  if rising_edge(clock_c) then
    if i5 = "1" then
      n27 <= "000000000000000000";
    elsif i4 = "1" then
      n27 <= n26;
    end if;
  end if;
end process;
n28 <= n24 + n27;
process (clock_c) begin
  if rising_edge(clock_c) then
    if i5 = "1" then
      n29 <= "000000000000000000";
    elsif i4 = "1" then
      n29 <= n28;
    end if;
  end if;
end process;
n30 <= n8 + n21;
n31 <= n10 + n29;
n32 <= n30 & n31;
process (clock_c) begin
  if rising_edge(clock_c) then
    if i5 = "1" then
      n33 <= "000000000000000000000000000000000000";
    elsif i4 = "1" then
      n33 <= n32;
    end if;
  end if;
end process;
n34 <= n8 - n21;
n35 <= n10 - n29;
n36 <= n34 & n35;
process (clock_c) begin
  if rising_edge(clock_c) then
    if i5 = "1" then
      n37 <= "000000000000000000000000000000000000";
    elsif i4 = "1" then
      n37 <= n36;
    end if;
  end if;
end process;
o2 <= n37;
o1 <= n33;
end architecture rtl;

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
entity cf_fft_256_18_4 is
port (
clock_c : in std_logic;
i1 : in  unsigned(0 downto 0);
i2 : in  unsigned(35 downto 0);
i3 : in  unsigned(35 downto 0);
i4 : in  unsigned(0 downto 0);
i5 : in  unsigned(0 downto 0);
o1 : out unsigned(0 downto 0);
o2 : out unsigned(35 downto 0);
o3 : out unsigned(35 downto 0));
end entity cf_fft_256_18_4;
architecture rtl of cf_fft_256_18_4 is
signal n1 : unsigned(0 downto 0);
signal n2 : unsigned(71 downto 0);
signal n3 : unsigned(0 downto 0) := "0";
signal n4 : unsigned(0 downto 0) := "0";
signal n5 : unsigned(0 downto 0) := "0";
signal n6 : unsigned(0 downto 0) := "0";
signal n7 : unsigned(5 downto 0);
signal n8 : unsigned(5 downto 0) := "000000";
signal n9 : unsigned(5 downto 0) := "000000";
signal n10 : unsigned(5 downto 0) := "000000";
signal n11 : unsigned(5 downto 0) := "000000";
signal n12 : unsigned(0 downto 0);
signal n13 : unsigned(0 downto 0) := "0";
signal n14 : unsigned(0 downto 0) := "0";
signal n15 : unsigned(0 downto 0) := "0";
signal n16 : unsigned(0 downto 0) := "0";
signal n17 : unsigned(0 downto 0);
signal n18 : unsigned(1 downto 0);
signal n19 : unsigned(35 downto 0);
signal n20 : unsigned(35 downto 0);
signal n21 : unsigned(35 downto 0);
signal n22 : unsigned(35 downto 0);
signal n23 : unsigned(35 downto 0);
signal n24 : unsigned(35 downto 0);
signal s25_1 : unsigned(0 downto 0);
signal s26_1 : unsigned(35 downto 0);
signal s26_2 : unsigned(35 downto 0);
signal s27_1 : unsigned(6 downto 0);
signal s27_2 : unsigned(0 downto 0);
signal s28_1 : unsigned(0 downto 0);
signal s28_2 : unsigned(0 downto 0);
signal s28_3 : unsigned(71 downto 0);
signal s29_1 : unsigned(71 downto 0);
component cf_fft_256_18_30 is
port (
clock_c : in std_logic;
i1 : in  unsigned(1 downto 0);
i2 : in  unsigned(0 downto 0);
i3 : in  unsigned(0 downto 0);
o1 : out unsigned(0 downto 0));
end component cf_fft_256_18_30;
component cf_fft_256_18_5 is
port (
clock_c : in std_logic;
i1 : in  unsigned(35 downto 0);
i2 : in  unsigned(35 downto 0);
i3 : in  unsigned(0 downto 0);
i4 : in  unsigned(0 downto 0);
i5 : in  unsigned(0 downto 0);
o1 : out unsigned(35 downto 0);
o2 : out unsigned(35 downto 0));
end component cf_fft_256_18_5;
component cf_fft_256_18_21 is
port (
clock_c : in std_logic;
i1 : in  unsigned(0 downto 0);
i2 : in  unsigned(0 downto 0);
i3 : in  unsigned(0 downto 0);
o1 : out unsigned(6 downto 0);
o2 : out unsigned(0 downto 0));
end component cf_fft_256_18_21;
component cf_fft_256_18_18 is
port (
clock_c : in std_logic;
i1 : in  unsigned(71 downto 0);
i2 : in  unsigned(0 downto 0);
i3 : in  unsigned(5 downto 0);
i4 : in  unsigned(0 downto 0);
i5 : in  unsigned(0 downto 0);
i6 : in  unsigned(0 downto 0);
o1 : out unsigned(0 downto 0);
o2 : out unsigned(0 downto 0);
o3 : out unsigned(71 downto 0));
end component cf_fft_256_18_18;
component cf_fft_256_18_17 is
port (
clock_c : in std_logic;
i1 : in  unsigned(71 downto 0);
i2 : in  unsigned(0 downto 0);
i3 : in  unsigned(5 downto 0);
i4 : in  unsigned(0 downto 0);
i5 : in  unsigned(0 downto 0);
i6 : in  unsigned(0 downto 0);
o1 : out unsigned(71 downto 0));
end component cf_fft_256_18_17;
begin
n1 <= s27_1(6 downto 6);
n2 <= s26_1 & s26_2;
process (clock_c) begin
  if rising_edge(clock_c) then
    if i5 = "1" then
      n3 <= "0";
    elsif i4 = "1" then
      n3 <= s27_2;
    end if;
  end if;
end process;
process (clock_c) begin
  if rising_edge(clock_c) then
    if i5 = "1" then
      n4 <= "0";
    elsif i4 = "1" then
      n4 <= n3;
    end if;
  end if;
end process;
process (clock_c) begin
  if rising_edge(clock_c) then
    if i5 = "1" then
      n5 <= "0";
    elsif i4 = "1" then
      n5 <= n4;
    end if;
  end if;
end process;
process (clock_c) begin
  if rising_edge(clock_c) then
    if i5 = "1" then
      n6 <= "0";
    elsif i4 = "1" then
      n6 <= n5;
    end if;
  end if;
end process;
n7 <= s27_1(6 downto 6) &
  s27_1(5 downto 5) &
  s27_1(4 downto 4) &
  s27_1(3 downto 3) &
  s27_1(2 downto 2) &
  s27_1(1 downto 1);
process (clock_c) begin
  if rising_edge(clock_c) then
    if i5 = "1" then
      n8 <= "000000";
    elsif i4 = "1" then
      n8 <= n7;
    end if;
  end if;
end process;
process (clock_c) begin
  if rising_edge(clock_c) then
    if i5 = "1" then
      n9 <= "000000";
    elsif i4 = "1" then
      n9 <= n8;
    end if;
  end if;
end process;
process (clock_c) begin
  if rising_edge(clock_c) then
    if i5 = "1" then
      n10 <= "000000";
    elsif i4 = "1" then
      n10 <= n9;
    end if;
  end if;
end process;
process (clock_c) begin
  if rising_edge(clock_c) then
    if i5 = "1" then
      n11 <= "000000";
    elsif i4 = "1" then
      n11 <= n10;
    end if;
  end if;
end process;
n12 <= s27_1(0 downto 0);
process (clock_c) begin
  if rising_edge(clock_c) then
    if i5 = "1" then
      n13 <= "0";
    elsif i4 = "1" then
      n13 <= n12;
    end if;
  end if;
end process;
process (clock_c) begin
  if rising_edge(clock_c) then
    if i5 = "1" then
      n14 <= "0";
    elsif i4 = "1" then
      n14 <= n13;
    end if;
  end if;
end process;
process (clock_c) begin
  if rising_edge(clock_c) then
    if i5 = "1" then
      n15 <= "0";
    elsif i4 = "1" then
      n15 <= n14;
    end if;
  end if;
end process;
process (clock_c) begin
  if rising_edge(clock_c) then
    if i5 = "1" then
      n16 <= "0";
    elsif i4 = "1" then
      n16 <= n15;
    end if;
  end if;
end process;
n17 <= not n16;
n18 <= s28_2 & s28_1;
n19 <= s28_3(71 downto 71) &
  s28_3(70 downto 70) &
  s28_3(69 downto 69) &
  s28_3(68 downto 68) &
  s28_3(67 downto 67) &
  s28_3(66 downto 66) &
  s28_3(65 downto 65) &
  s28_3(64 downto 64) &
  s28_3(63 downto 63) &
  s28_3(62 downto 62) &
  s28_3(61 downto 61) &
  s28_3(60 downto 60) &
  s28_3(59 downto 59) &
  s28_3(58 downto 58) &
  s28_3(57 downto 57) &
  s28_3(56 downto 56) &
  s28_3(55 downto 55) &
  s28_3(54 downto 54) &
  s28_3(53 downto 53) &
  s28_3(52 downto 52) &
  s28_3(51 downto 51) &
  s28_3(50 downto 50) &
  s28_3(49 downto 49) &
  s28_3(48 downto 48) &
  s28_3(47 downto 47) &
  s28_3(46 downto 46) &
  s28_3(45 downto 45) &
  s28_3(44 downto 44) &
  s28_3(43 downto 43) &
  s28_3(42 downto 42) &
  s28_3(41 downto 41) &
  s28_3(40 downto 40) &
  s28_3(39 downto 39) &
  s28_3(38 downto 38) &
  s28_3(37 downto 37) &
  s28_3(36 downto 36);
n20 <= s28_3(35 downto 35) &
  s28_3(34 downto 34) &
  s28_3(33 downto 33) &
  s28_3(32 downto 32) &
  s28_3(31 downto 31) &
  s28_3(30 downto 30) &
  s28_3(29 downto 29) &
  s28_3(28 downto 28) &
  s28_3(27 downto 27) &
  s28_3(26 downto 26) &
  s28_3(25 downto 25) &
  s28_3(24 downto 24) &
  s28_3(23 downto 23) &
  s28_3(22 downto 22) &
  s28_3(21 downto 21) &
  s28_3(20 downto 20) &
  s28_3(19 downto 19) &
  s28_3(18 downto 18) &
  s28_3(17 downto 17) &
  s28_3(16 downto 16) &
  s28_3(15 downto 15) &
  s28_3(14 downto 14) &
  s28_3(13 downto 13) &
  s28_3(12 downto 12) &
  s28_3(11 downto 11) &
  s28_3(10 downto 10) &
  s28_3(9 downto 9) &
  s28_3(8 downto 8) &
  s28_3(7 downto 7) &
  s28_3(6 downto 6) &
  s28_3(5 downto 5) &
  s28_3(4 downto 4) &
  s28_3(3 downto 3) &
  s28_3(2 downto 2) &
  s28_3(1 downto 1) &
  s28_3(0 downto 0);
n21 <= s29_1(71 downto 71) &
  s29_1(70 downto 70) &
  s29_1(69 downto 69) &
  s29_1(68 downto 68) &
  s29_1(67 downto 67) &
  s29_1(66 downto 66) &
  s29_1(65 downto 65) &
  s29_1(64 downto 64) &
  s29_1(63 downto 63) &
  s29_1(62 downto 62) &
  s29_1(61 downto 61) &
  s29_1(60 downto 60) &
  s29_1(59 downto 59) &
  s29_1(58 downto 58) &
  s29_1(57 downto 57) &
  s29_1(56 downto 56) &
  s29_1(55 downto 55) &
  s29_1(54 downto 54) &
  s29_1(53 downto 53) &
  s29_1(52 downto 52) &
  s29_1(51 downto 51) &
  s29_1(50 downto 50) &
  s29_1(49 downto 49) &
  s29_1(48 downto 48) &
  s29_1(47 downto 47) &
  s29_1(46 downto 46) &
  s29_1(45 downto 45) &
  s29_1(44 downto 44) &
  s29_1(43 downto 43) &
  s29_1(42 downto 42) &
  s29_1(41 downto 41) &
  s29_1(40 downto 40) &
  s29_1(39 downto 39) &
  s29_1(38 downto 38) &
  s29_1(37 downto 37) &
  s29_1(36 downto 36);
n22 <= s29_1(35 downto 35) &
  s29_1(34 downto 34) &
  s29_1(33 downto 33) &
  s29_1(32 downto 32) &
  s29_1(31 downto 31) &
  s29_1(30 downto 30) &
  s29_1(29 downto 29) &
  s29_1(28 downto 28) &
  s29_1(27 downto 27) &
  s29_1(26 downto 26) &
  s29_1(25 downto 25) &
  s29_1(24 downto 24) &
  s29_1(23 downto 23) &
  s29_1(22 downto 22) &
  s29_1(21 downto 21) &
  s29_1(20 downto 20) &
  s29_1(19 downto 19) &
  s29_1(18 downto 18) &
  s29_1(17 downto 17) &
  s29_1(16 downto 16) &
  s29_1(15 downto 15) &
  s29_1(14 downto 14) &
  s29_1(13 downto 13) &
  s29_1(12 downto 12) &
  s29_1(11 downto 11) &
  s29_1(10 downto 10) &
  s29_1(9 downto 9) &
  s29_1(8 downto 8) &
  s29_1(7 downto 7) &
  s29_1(6 downto 6) &
  s29_1(5 downto 5) &
  s29_1(4 downto 4) &
  s29_1(3 downto 3) &
  s29_1(2 downto 2) &
  s29_1(1 downto 1) &
  s29_1(0 downto 0);
n23 <= n20 when s25_1 = "1" else n19;
n24 <= n22 when s25_1 = "1" else n21;
s25 : cf_fft_256_18_30 port map (clock_c, n18, i4, i5, s25_1);
s26 : cf_fft_256_18_5 port map (clock_c, i2, i3, n1, i4, i5, s26_1, s26_2);
s27 : cf_fft_256_18_21 port map (clock_c, i1, i4, i5, s27_1, s27_2);
s28 : cf_fft_256_18_18 port map (clock_c, n2, n6, n11, n17, i4, i5, s28_1, s28_2, s28_3);
s29 : cf_fft_256_18_17 port map (clock_c, n2, n6, n11, n16, i4, i5, s29_1);
o3 <= n24;
o2 <= n23;
o1 <= s28_1;
end architecture rtl;

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
entity cf_fft_256_18_3 is
port (
clock_c : in std_logic;
i1 : in  unsigned(0 downto 0);
i2 : in  unsigned(35 downto 0);
i3 : in  unsigned(35 downto 0);
i4 : in  unsigned(0 downto 0);
i5 : in  unsigned(0 downto 0);
o1 : out unsigned(0 downto 0);
o2 : out unsigned(35 downto 0);
o3 : out unsigned(35 downto 0));
end entity cf_fft_256_18_3;
architecture rtl of cf_fft_256_18_3 is
signal n1 : unsigned(0 downto 0);
signal n2 : unsigned(71 downto 0);
signal n3 : unsigned(0 downto 0) := "0";
signal n4 : unsigned(0 downto 0) := "0";
signal n5 : unsigned(0 downto 0) := "0";
signal n6 : unsigned(0 downto 0) := "0";
signal n7 : unsigned(5 downto 0);
signal n8 : unsigned(5 downto 0) := "000000";
signal n9 : unsigned(5 downto 0) := "000000";
signal n10 : unsigned(5 downto 0) := "000000";
signal n11 : unsigned(5 downto 0) := "000000";
signal n12 : unsigned(0 downto 0);
signal n13 : unsigned(0 downto 0) := "0";
signal n14 : unsigned(0 downto 0) := "0";
signal n15 : unsigned(0 downto 0) := "0";
signal n16 : unsigned(0 downto 0) := "0";
signal n17 : unsigned(0 downto 0);
signal n18 : unsigned(1 downto 0);
signal n19 : unsigned(35 downto 0);
signal n20 : unsigned(35 downto 0);
signal n21 : unsigned(35 downto 0);
signal n22 : unsigned(35 downto 0);
signal n23 : unsigned(35 downto 0);
signal n24 : unsigned(35 downto 0);
signal s25_1 : unsigned(35 downto 0);
signal s25_2 : unsigned(35 downto 0);
signal s26_1 : unsigned(0 downto 0);
signal s27_1 : unsigned(0 downto 0);
signal s27_2 : unsigned(0 downto 0);
signal s27_3 : unsigned(71 downto 0);
signal s28_1 : unsigned(71 downto 0);
signal s29_1 : unsigned(6 downto 0);
signal s29_2 : unsigned(0 downto 0);
component cf_fft_256_18_5 is
port (
clock_c : in std_logic;
i1 : in  unsigned(35 downto 0);
i2 : in  unsigned(35 downto 0);
i3 : in  unsigned(0 downto 0);
i4 : in  unsigned(0 downto 0);
i5 : in  unsigned(0 downto 0);
o1 : out unsigned(35 downto 0);
o2 : out unsigned(35 downto 0));
end component cf_fft_256_18_5;
component cf_fft_256_18_30 is
port (
clock_c : in std_logic;
i1 : in  unsigned(1 downto 0);
i2 : in  unsigned(0 downto 0);
i3 : in  unsigned(0 downto 0);
o1 : out unsigned(0 downto 0));
end component cf_fft_256_18_30;
component cf_fft_256_18_18 is
port (
clock_c : in std_logic;
i1 : in  unsigned(71 downto 0);
i2 : in  unsigned(0 downto 0);
i3 : in  unsigned(5 downto 0);
i4 : in  unsigned(0 downto 0);
i5 : in  unsigned(0 downto 0);
i6 : in  unsigned(0 downto 0);
o1 : out unsigned(0 downto 0);
o2 : out unsigned(0 downto 0);
o3 : out unsigned(71 downto 0));
end component cf_fft_256_18_18;
component cf_fft_256_18_17 is
port (
clock_c : in std_logic;
i1 : in  unsigned(71 downto 0);
i2 : in  unsigned(0 downto 0);
i3 : in  unsigned(5 downto 0);
i4 : in  unsigned(0 downto 0);
i5 : in  unsigned(0 downto 0);
i6 : in  unsigned(0 downto 0);
o1 : out unsigned(71 downto 0));
end component cf_fft_256_18_17;
component cf_fft_256_18_21 is
port (
clock_c : in std_logic;
i1 : in  unsigned(0 downto 0);
i2 : in  unsigned(0 downto 0);
i3 : in  unsigned(0 downto 0);
o1 : out unsigned(6 downto 0);
o2 : out unsigned(0 downto 0));
end component cf_fft_256_18_21;
begin
n1 <= "0";
n2 <= s25_1 & s25_2;
process (clock_c) begin
  if rising_edge(clock_c) then
    if i5 = "1" then
      n3 <= "0";
    elsif i4 = "1" then
      n3 <= s29_2;
    end if;
  end if;
end process;
process (clock_c) begin
  if rising_edge(clock_c) then
    if i5 = "1" then
      n4 <= "0";
    elsif i4 = "1" then
      n4 <= n3;
    end if;
  end if;
end process;
process (clock_c) begin
  if rising_edge(clock_c) then
    if i5 = "1" then
      n5 <= "0";
    elsif i4 = "1" then
      n5 <= n4;
    end if;
  end if;
end process;
process (clock_c) begin
  if rising_edge(clock_c) then
    if i5 = "1" then
      n6 <= "0";
    elsif i4 = "1" then
      n6 <= n5;
    end if;
  end if;
end process;
n7 <= s29_1(6 downto 6) &
  s29_1(5 downto 5) &
  s29_1(4 downto 4) &
  s29_1(3 downto 3) &
  s29_1(2 downto 2) &
  s29_1(1 downto 1);
process (clock_c) begin
  if rising_edge(clock_c) then
    if i5 = "1" then
      n8 <= "000000";
    elsif i4 = "1" then
      n8 <= n7;
    end if;
  end if;
end process;
process (clock_c) begin
  if rising_edge(clock_c) then
    if i5 = "1" then
      n9 <= "000000";
    elsif i4 = "1" then
      n9 <= n8;
    end if;
  end if;
end process;
process (clock_c) begin
  if rising_edge(clock_c) then
    if i5 = "1" then
      n10 <= "000000";
    elsif i4 = "1" then
      n10 <= n9;
    end if;
  end if;
end process;
process (clock_c) begin
  if rising_edge(clock_c) then
    if i5 = "1" then
      n11 <= "000000";
    elsif i4 = "1" then
      n11 <= n10;
    end if;
  end if;
end process;
n12 <= s29_1(0 downto 0);
process (clock_c) begin
  if rising_edge(clock_c) then
    if i5 = "1" then
      n13 <= "0";
    elsif i4 = "1" then
      n13 <= n12;
    end if;
  end if;
end process;
process (clock_c) begin
  if rising_edge(clock_c) then
    if i5 = "1" then
      n14 <= "0";
    elsif i4 = "1" then
      n14 <= n13;
    end if;
  end if;
end process;
process (clock_c) begin
  if rising_edge(clock_c) then
    if i5 = "1" then
      n15 <= "0";
    elsif i4 = "1" then
      n15 <= n14;
    end if;
  end if;
end process;
process (clock_c) begin
  if rising_edge(clock_c) then
    if i5 = "1" then
      n16 <= "0";
    elsif i4 = "1" then
      n16 <= n15;
    end if;
  end if;
end process;
n17 <= not n16;
n18 <= s27_2 & s27_1;
n19 <= s27_3(71 downto 71) &
  s27_3(70 downto 70) &
  s27_3(69 downto 69) &
  s27_3(68 downto 68) &
  s27_3(67 downto 67) &
  s27_3(66 downto 66) &
  s27_3(65 downto 65) &
  s27_3(64 downto 64) &
  s27_3(63 downto 63) &
  s27_3(62 downto 62) &
  s27_3(61 downto 61) &
  s27_3(60 downto 60) &
  s27_3(59 downto 59) &
  s27_3(58 downto 58) &
  s27_3(57 downto 57) &
  s27_3(56 downto 56) &
  s27_3(55 downto 55) &
  s27_3(54 downto 54) &
  s27_3(53 downto 53) &
  s27_3(52 downto 52) &
  s27_3(51 downto 51) &
  s27_3(50 downto 50) &
  s27_3(49 downto 49) &
  s27_3(48 downto 48) &
  s27_3(47 downto 47) &
  s27_3(46 downto 46) &
  s27_3(45 downto 45) &
  s27_3(44 downto 44) &
  s27_3(43 downto 43) &
  s27_3(42 downto 42) &
  s27_3(41 downto 41) &
  s27_3(40 downto 40) &
  s27_3(39 downto 39) &
  s27_3(38 downto 38) &
  s27_3(37 downto 37) &
  s27_3(36 downto 36);
n20 <= s27_3(35 downto 35) &
  s27_3(34 downto 34) &
  s27_3(33 downto 33) &
  s27_3(32 downto 32) &
  s27_3(31 downto 31) &
  s27_3(30 downto 30) &
  s27_3(29 downto 29) &
  s27_3(28 downto 28) &
  s27_3(27 downto 27) &
  s27_3(26 downto 26) &
  s27_3(25 downto 25) &
  s27_3(24 downto 24) &
  s27_3(23 downto 23) &
  s27_3(22 downto 22) &
  s27_3(21 downto 21) &
  s27_3(20 downto 20) &
  s27_3(19 downto 19) &
  s27_3(18 downto 18) &
  s27_3(17 downto 17) &
  s27_3(16 downto 16) &
  s27_3(15 downto 15) &
  s27_3(14 downto 14) &
  s27_3(13 downto 13) &
  s27_3(12 downto 12) &
  s27_3(11 downto 11) &
  s27_3(10 downto 10) &
  s27_3(9 downto 9) &
  s27_3(8 downto 8) &
  s27_3(7 downto 7) &
  s27_3(6 downto 6) &
  s27_3(5 downto 5) &
  s27_3(4 downto 4) &
  s27_3(3 downto 3) &
  s27_3(2 downto 2) &
  s27_3(1 downto 1) &
  s27_3(0 downto 0);
n21 <= s28_1(71 downto 71) &
  s28_1(70 downto 70) &
  s28_1(69 downto 69) &
  s28_1(68 downto 68) &
  s28_1(67 downto 67) &
  s28_1(66 downto 66) &
  s28_1(65 downto 65) &
  s28_1(64 downto 64) &
  s28_1(63 downto 63) &
  s28_1(62 downto 62) &
  s28_1(61 downto 61) &
  s28_1(60 downto 60) &
  s28_1(59 downto 59) &
  s28_1(58 downto 58) &
  s28_1(57 downto 57) &
  s28_1(56 downto 56) &
  s28_1(55 downto 55) &
  s28_1(54 downto 54) &
  s28_1(53 downto 53) &
  s28_1(52 downto 52) &
  s28_1(51 downto 51) &
  s28_1(50 downto 50) &
  s28_1(49 downto 49) &
  s28_1(48 downto 48) &
  s28_1(47 downto 47) &
  s28_1(46 downto 46) &
  s28_1(45 downto 45) &
  s28_1(44 downto 44) &
  s28_1(43 downto 43) &
  s28_1(42 downto 42) &
  s28_1(41 downto 41) &
  s28_1(40 downto 40) &
  s28_1(39 downto 39) &
  s28_1(38 downto 38) &
  s28_1(37 downto 37) &
  s28_1(36 downto 36);
n22 <= s28_1(35 downto 35) &
  s28_1(34 downto 34) &
  s28_1(33 downto 33) &
  s28_1(32 downto 32) &
  s28_1(31 downto 31) &
  s28_1(30 downto 30) &
  s28_1(29 downto 29) &
  s28_1(28 downto 28) &
  s28_1(27 downto 27) &
  s28_1(26 downto 26) &
  s28_1(25 downto 25) &
  s28_1(24 downto 24) &
  s28_1(23 downto 23) &
  s28_1(22 downto 22) &
  s28_1(21 downto 21) &
  s28_1(20 downto 20) &
  s28_1(19 downto 19) &
  s28_1(18 downto 18) &
  s28_1(17 downto 17) &
  s28_1(16 downto 16) &
  s28_1(15 downto 15) &
  s28_1(14 downto 14) &
  s28_1(13 downto 13) &
  s28_1(12 downto 12) &
  s28_1(11 downto 11) &
  s28_1(10 downto 10) &
  s28_1(9 downto 9) &
  s28_1(8 downto 8) &
  s28_1(7 downto 7) &
  s28_1(6 downto 6) &
  s28_1(5 downto 5) &
  s28_1(4 downto 4) &
  s28_1(3 downto 3) &
  s28_1(2 downto 2) &
  s28_1(1 downto 1) &
  s28_1(0 downto 0);
n23 <= n20 when s26_1 = "1" else n19;
n24 <= n22 when s26_1 = "1" else n21;
s25 : cf_fft_256_18_5 port map (clock_c, i2, i3, n1, i4, i5, s25_1, s25_2);
s26 : cf_fft_256_18_30 port map (clock_c, n18, i4, i5, s26_1);
s27 : cf_fft_256_18_18 port map (clock_c, n2, n6, n11, n17, i4, i5, s27_1, s27_2, s27_3);
s28 : cf_fft_256_18_17 port map (clock_c, n2, n6, n11, n16, i4, i5, s28_1);
s29 : cf_fft_256_18_21 port map (clock_c, i1, i4, i5, s29_1, s29_2);
o3 <= n24;
o2 <= n23;
o1 <= s27_1;
end architecture rtl;

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
entity cf_fft_256_18_2 is
port (
clock_c : in std_logic;
i1 : in  unsigned(0 downto 0);
i2 : in  unsigned(35 downto 0);
i3 : in  unsigned(35 downto 0);
i4 : in  unsigned(0 downto 0);
i5 : in  unsigned(0 downto 0);
o1 : out unsigned(0 downto 0);
o2 : out unsigned(35 downto 0);
o3 : out unsigned(35 downto 0));
end entity cf_fft_256_18_2;
architecture rtl of cf_fft_256_18_2 is
signal s1_1 : unsigned(0 downto 0);
signal s1_2 : unsigned(35 downto 0);
signal s1_3 : unsigned(35 downto 0);
signal s2_1 : unsigned(0 downto 0);
signal s2_2 : unsigned(35 downto 0);
signal s2_3 : unsigned(35 downto 0);
signal s3_1 : unsigned(0 downto 0);
signal s3_2 : unsigned(35 downto 0);
signal s3_3 : unsigned(35 downto 0);
signal s4_1 : unsigned(0 downto 0);
signal s4_2 : unsigned(35 downto 0);
signal s4_3 : unsigned(35 downto 0);
signal s5_1 : unsigned(0 downto 0);
signal s5_2 : unsigned(35 downto 0);
signal s5_3 : unsigned(35 downto 0);
signal s6_1 : unsigned(0 downto 0);
signal s6_2 : unsigned(35 downto 0);
signal s6_3 : unsigned(35 downto 0);
signal s7_1 : unsigned(0 downto 0);
signal s7_2 : unsigned(35 downto 0);
signal s7_3 : unsigned(35 downto 0);
signal s8_1 : unsigned(0 downto 0);
signal s8_2 : unsigned(35 downto 0);
signal s8_3 : unsigned(35 downto 0);
component cf_fft_256_18_16 is
port (
clock_c : in std_logic;
i1 : in  unsigned(0 downto 0);
i2 : in  unsigned(35 downto 0);
i3 : in  unsigned(35 downto 0);
i4 : in  unsigned(0 downto 0);
i5 : in  unsigned(0 downto 0);
o1 : out unsigned(0 downto 0);
o2 : out unsigned(35 downto 0);
o3 : out unsigned(35 downto 0));
end component cf_fft_256_18_16;
component cf_fft_256_18_14 is
port (
clock_c : in std_logic;
i1 : in  unsigned(0 downto 0);
i2 : in  unsigned(35 downto 0);
i3 : in  unsigned(35 downto 0);
i4 : in  unsigned(0 downto 0);
i5 : in  unsigned(0 downto 0);
o1 : out unsigned(0 downto 0);
o2 : out unsigned(35 downto 0);
o3 : out unsigned(35 downto 0));
end component cf_fft_256_18_14;
component cf_fft_256_18_12 is
port (
clock_c : in std_logic;
i1 : in  unsigned(0 downto 0);
i2 : in  unsigned(35 downto 0);
i3 : in  unsigned(35 downto 0);
i4 : in  unsigned(0 downto 0);
i5 : in  unsigned(0 downto 0);
o1 : out unsigned(0 downto 0);
o2 : out unsigned(35 downto 0);
o3 : out unsigned(35 downto 0));
end component cf_fft_256_18_12;
component cf_fft_256_18_10 is
port (
clock_c : in std_logic;
i1 : in  unsigned(0 downto 0);
i2 : in  unsigned(35 downto 0);
i3 : in  unsigned(35 downto 0);
i4 : in  unsigned(0 downto 0);
i5 : in  unsigned(0 downto 0);
o1 : out unsigned(0 downto 0);
o2 : out unsigned(35 downto 0);
o3 : out unsigned(35 downto 0));
end component cf_fft_256_18_10;
component cf_fft_256_18_8 is
port (
clock_c : in std_logic;
i1 : in  unsigned(0 downto 0);
i2 : in  unsigned(35 downto 0);
i3 : in  unsigned(35 downto 0);
i4 : in  unsigned(0 downto 0);
i5 : in  unsigned(0 downto 0);
o1 : out unsigned(0 downto 0);
o2 : out unsigned(35 downto 0);
o3 : out unsigned(35 downto 0));
end component cf_fft_256_18_8;
component cf_fft_256_18_6 is
port (
clock_c : in std_logic;
i1 : in  unsigned(0 downto 0);
i2 : in  unsigned(35 downto 0);
i3 : in  unsigned(35 downto 0);
i4 : in  unsigned(0 downto 0);
i5 : in  unsigned(0 downto 0);
o1 : out unsigned(0 downto 0);
o2 : out unsigned(35 downto 0);
o3 : out unsigned(35 downto 0));
end component cf_fft_256_18_6;
component cf_fft_256_18_4 is
port (
clock_c : in std_logic;
i1 : in  unsigned(0 downto 0);
i2 : in  unsigned(35 downto 0);
i3 : in  unsigned(35 downto 0);
i4 : in  unsigned(0 downto 0);
i5 : in  unsigned(0 downto 0);
o1 : out unsigned(0 downto 0);
o2 : out unsigned(35 downto 0);
o3 : out unsigned(35 downto 0));
end component cf_fft_256_18_4;
component cf_fft_256_18_3 is
port (
clock_c : in std_logic;
i1 : in  unsigned(0 downto 0);
i2 : in  unsigned(35 downto 0);
i3 : in  unsigned(35 downto 0);
i4 : in  unsigned(0 downto 0);
i5 : in  unsigned(0 downto 0);
o1 : out unsigned(0 downto 0);
o2 : out unsigned(35 downto 0);
o3 : out unsigned(35 downto 0));
end component cf_fft_256_18_3;
begin
s1 : cf_fft_256_18_16 port map (clock_c, s3_1, s3_2, s3_3, i4, i5, s1_1, s1_2, s1_3);
s2 : cf_fft_256_18_14 port map (clock_c, s1_1, s1_2, s1_3, i4, i5, s2_1, s2_2, s2_3);
s3 : cf_fft_256_18_12 port map (clock_c, s4_1, s4_2, s4_3, i4, i5, s3_1, s3_2, s3_3);
s4 : cf_fft_256_18_10 port map (clock_c, s5_1, s5_2, s5_3, i4, i5, s4_1, s4_2, s4_3);
s5 : cf_fft_256_18_8 port map (clock_c, s6_1, s6_2, s6_3, i4, i5, s5_1, s5_2, s5_3);
s6 : cf_fft_256_18_6 port map (clock_c, s7_1, s7_2, s7_3, i4, i5, s6_1, s6_2, s6_3);
s7 : cf_fft_256_18_4 port map (clock_c, s8_1, s8_2, s8_3, i4, i5, s7_1, s7_2, s7_3);
s8 : cf_fft_256_18_3 port map (clock_c, i1, i2, i3, i4, i5, s8_1, s8_2, s8_3);
o3 <= s2_3;
o2 <= s2_2;
o1 <= s2_1;
end architecture rtl;

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
entity cf_fft_256_18_1 is
port (
clock_c : in std_logic;
i1 : in  unsigned(0 downto 0);
i2 : in  unsigned(35 downto 0);
i3 : in  unsigned(35 downto 0);
i4 : in  unsigned(0 downto 0);
i5 : in  unsigned(0 downto 0);
o1 : out unsigned(0 downto 0);
o2 : out unsigned(35 downto 0);
o3 : out unsigned(35 downto 0));
end entity cf_fft_256_18_1;
architecture rtl of cf_fft_256_18_1 is
signal s1_1 : unsigned(0 downto 0);
signal s1_2 : unsigned(35 downto 0);
signal s1_3 : unsigned(35 downto 0);
signal s2_1 : unsigned(0 downto 0);
signal s2_2 : unsigned(35 downto 0);
signal s2_3 : unsigned(35 downto 0);
component cf_fft_256_18_20 is
port (
clock_c : in std_logic;
i1 : in  unsigned(0 downto 0);
i2 : in  unsigned(35 downto 0);
i3 : in  unsigned(35 downto 0);
i4 : in  unsigned(0 downto 0);
i5 : in  unsigned(0 downto 0);
o1 : out unsigned(0 downto 0);
o2 : out unsigned(35 downto 0);
o3 : out unsigned(35 downto 0));
end component cf_fft_256_18_20;
component cf_fft_256_18_2 is
port (
clock_c : in std_logic;
i1 : in  unsigned(0 downto 0);
i2 : in  unsigned(35 downto 0);
i3 : in  unsigned(35 downto 0);
i4 : in  unsigned(0 downto 0);
i5 : in  unsigned(0 downto 0);
o1 : out unsigned(0 downto 0);
o2 : out unsigned(35 downto 0);
o3 : out unsigned(35 downto 0));
end component cf_fft_256_18_2;
begin
s1 : cf_fft_256_18_20 port map (clock_c, i1, i2, i3, i4, i5, s1_1, s1_2, s1_3);
s2 : cf_fft_256_18_2 port map (clock_c, s1_1, s1_2, s1_3, i4, i5, s2_1, s2_2, s2_3);
o3 <= s2_3;
o2 <= s2_2;
o1 <= s2_1;
end architecture rtl;

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
entity cf_fft_256_18 is
port(
signal clock_c : in std_logic;
signal enable_i : in unsigned(0 downto 0);
signal reset_i : in unsigned(0 downto 0);
signal sync_i : in unsigned(0 downto 0);
signal data_0_i : in unsigned(35 downto 0);
signal data_1_i : in unsigned(35 downto 0);
signal sync_o : out unsigned(0 downto 0);
signal data_0_o : out unsigned(35 downto 0);
signal data_1_o : out unsigned(35 downto 0));
end entity cf_fft_256_18;
architecture rtl of cf_fft_256_18 is
component cf_fft_256_18_1 is
port (
clock_c : in std_logic;
i1 : in  unsigned(0 downto 0);
i2 : in  unsigned(35 downto 0);
i3 : in  unsigned(35 downto 0);
i4 : in  unsigned(0 downto 0);
i5 : in  unsigned(0 downto 0);
o1 : out unsigned(0 downto 0);
o2 : out unsigned(35 downto 0);
o3 : out unsigned(35 downto 0));
end component cf_fft_256_18_1;
signal n1 : unsigned(0 downto 0);
signal n2 : unsigned(35 downto 0);
signal n3 : unsigned(35 downto 0);
begin
s1 : cf_fft_256_18_1 port map (clock_c, sync_i, data_0_i, data_1_i, enable_i, reset_i, n1, n2, n3);
sync_o <= n1;
data_0_o <= n2;
data_1_o <= n3;
end architecture rtl;


