--
--  Copyright (c) 2003 Launchbird Design Systems, Inc.
--  All rights reserved.
--  
--  Redistribution and use in source and binary forms, with or without modification, are permitted provided that the following conditions are met:
--    Redistributions of source code must retain the above copyright notice, this list of conditions and the following disclaimer.
--    Redistributions in binary form must reproduce the above copyright notice, this list of conditions and the following disclaimer in the documentation and/or other materials provided with the distribution.
--  
--  THIS SOFTWARE IS PROVIDED BY THE COPYRIGHT HOLDERS AND CONTRIBUTORS "AS IS" AND ANY EXPRESS OR IMPLIED WARRANTIES,
--  INCLUDING, BUT NOT LIMITED TO, THE IMPLIED WARRANTIES OF MERCHANTABILITY AND FITNESS FOR A PARTICULAR PURPOSE ARE DISCLAIMED.
--  IN NO EVENT SHALL THE COPYRIGHT OWNER OR CONTRIBUTORS BE LIABLE FOR ANY DIRECT, INDIRECT, INCIDENTAL, SPECIAL, EXEMPLARY,
--  OR CONSEQUENTIAL DAMAGES (INCLUDING, BUT NOT LIMITED TO, PROCUREMENT OF SUBSTITUTE GOODS OR SERVICES; LOSS OF USE, DATA, OR PROFITS;
--  OR BUSINESS INTERRUPTION) HOWEVER CAUSED AND ON ANY THEORY OF LIABILITY, WHETHER IN CONTRACT, STRICT LIABILITY, OR TORT
--  (INCLUDING NEGLIGENCE OR OTHERWISE) ARISING IN ANY WAY OUT OF THE USE OF THIS SOFTWARE, EVEN IF ADVISED OF THE POSSIBILITY OF SUCH DAMAGE.
--  
--  
--  Overview:
--  
--    Performs a radix 2 Fast Fourier Transform.
--    The FFT architecture is pipelined on a rank basis; each rank has its own butterfly and ranks are
--    isolated from each other using memory interleavers.  This FFT can perform calcualations on continuous
--    streaming data (one data set right after another).  More over, inputs and outputs are passed in pairs,
--    doubling the bandwidth.  For instance, a 2048 point FFT can perform a transform every 1024 cycles.
--  
--  Interface:
--  
--    Synchronization:
--      clock_c  : Clock input.
--      enable_i : Synchronous enable.
--      reset_i  : Synchronous reset.
--  
--    Inputs:
--      sync_i     : Input sync pulse must occur one frame prior to data input.
--      data_0_i   : Input data 0.  Width is 2 * precision.  Real on the left, imag on the right.
--      data_1_i   : Input data 1.  Width is 2 * precision.  Real on the left, imag on the right.
--  
--    Outputs:
--      sync_o     : Output sync pulse occurs one frame before data output.
--      data_0_o   : Output data 0.  Width is 2 * precision.  Real on the left, imag on the right.
--      data_1_o   : Output data 1.  Width is 2 * precision.  Real on the left, imag on the right.
--  
--  Built In Parameters:
--  
--    FFT Points   = 2048
--    Precision    = 16
--  
--  
--  
--  
--  Generated by Confluence 0.6.3  --  Launchbird Design Systems, Inc.  --  www.launchbird.com
--  
--  Build Date : Fri Aug 22 08:44:21 CDT 2003
--  
--  Interface
--  
--    Build Name    : cf_fft_2048_16
--    Clock Domains : clock_c  
--    Vector Input  : enable_i(1)
--    Vector Input  : reset_i(1)
--    Vector Input  : sync_i(1)
--    Vector Input  : data_0_i(32)
--    Vector Input  : data_1_i(32)
--    Vector Output : sync_o(1)
--    Vector Output : data_0_o(32)
--    Vector Output : data_1_o(32)
--  
--  
--  

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
entity cf_fft_2048_16_41 is
port (
clock_c : in std_logic;
i1 : in  unsigned(31 downto 0);
i2 : in  unsigned(31 downto 0);
i3 : in  unsigned(1 downto 0);
i4 : in  unsigned(0 downto 0);
i5 : in  unsigned(0 downto 0);
o1 : out unsigned(31 downto 0);
o2 : out unsigned(31 downto 0));
end entity cf_fft_2048_16_41;
architecture rtl of cf_fft_2048_16_41 is
signal n1 : unsigned(31 downto 0) := "00000000000000000000000000000000";
signal n2 : unsigned(15 downto 0);
signal n3 : unsigned(15 downto 0);
signal n4 : unsigned(31 downto 0) := "00000000000000000000000000000000";
signal n5 : unsigned(15 downto 0);
signal n6 : unsigned(15 downto 0);
signal n7 : unsigned(15 downto 0) := "0000000000000000";
signal n8 : unsigned(15 downto 0) := "0000000000000000";
signal n9 : unsigned(15 downto 0) := "0000000000000000";
signal n10 : unsigned(15 downto 0) := "0000000000000000";
signal n11 : unsigned(31 downto 0) := "00000000000000000000000000000000";
signal n12 : unsigned(15 downto 0);
signal n13 : unsigned(15 downto 0);
signal n14 : unsigned(31 downto 0);
signal n15 : unsigned(15 downto 0);
signal n16 : unsigned(15 downto 0) := "0000000000000000";
signal n17 : unsigned(31 downto 0);
signal n18 : unsigned(15 downto 0);
signal n19 : unsigned(15 downto 0) := "0000000000000000";
signal n20 : unsigned(15 downto 0);
signal n21 : unsigned(15 downto 0) := "0000000000000000";
signal n22 : unsigned(31 downto 0);
signal n23 : unsigned(15 downto 0);
signal n24 : unsigned(15 downto 0) := "0000000000000000";
signal n25 : unsigned(31 downto 0);
signal n26 : unsigned(15 downto 0);
signal n27 : unsigned(15 downto 0) := "0000000000000000";
signal n28 : unsigned(15 downto 0);
signal n29 : unsigned(15 downto 0) := "0000000000000000";
signal n30 : unsigned(15 downto 0);
signal n31 : unsigned(15 downto 0);
signal n32 : unsigned(31 downto 0);
signal n33 : unsigned(31 downto 0) := "00000000000000000000000000000000";
signal n34 : unsigned(15 downto 0);
signal n35 : unsigned(15 downto 0);
signal n36 : unsigned(31 downto 0);
signal n37 : unsigned(31 downto 0) := "00000000000000000000000000000000";
begin
process (clock_c) begin
  if rising_edge(clock_c) then
    if i5 = "1" then
      n1 <= "00000000000000000000000000000000";
    elsif i4 = "1" then
      n1 <= i1;
    end if;
  end if;
end process;
n2 <= n1(31 downto 31) &
  n1(30 downto 30) &
  n1(29 downto 29) &
  n1(28 downto 28) &
  n1(27 downto 27) &
  n1(26 downto 26) &
  n1(25 downto 25) &
  n1(24 downto 24) &
  n1(23 downto 23) &
  n1(22 downto 22) &
  n1(21 downto 21) &
  n1(20 downto 20) &
  n1(19 downto 19) &
  n1(18 downto 18) &
  n1(17 downto 17) &
  n1(16 downto 16);
n3 <= n1(15 downto 15) &
  n1(14 downto 14) &
  n1(13 downto 13) &
  n1(12 downto 12) &
  n1(11 downto 11) &
  n1(10 downto 10) &
  n1(9 downto 9) &
  n1(8 downto 8) &
  n1(7 downto 7) &
  n1(6 downto 6) &
  n1(5 downto 5) &
  n1(4 downto 4) &
  n1(3 downto 3) &
  n1(2 downto 2) &
  n1(1 downto 1) &
  n1(0 downto 0);
process (clock_c) begin
  if rising_edge(clock_c) then
    if i5 = "1" then
      n4 <= "00000000000000000000000000000000";
    elsif i4 = "1" then
      n4 <= i2;
    end if;
  end if;
end process;
n5 <= n4(31 downto 31) &
  n4(30 downto 30) &
  n4(29 downto 29) &
  n4(28 downto 28) &
  n4(27 downto 27) &
  n4(26 downto 26) &
  n4(25 downto 25) &
  n4(24 downto 24) &
  n4(23 downto 23) &
  n4(22 downto 22) &
  n4(21 downto 21) &
  n4(20 downto 20) &
  n4(19 downto 19) &
  n4(18 downto 18) &
  n4(17 downto 17) &
  n4(16 downto 16);
n6 <= n4(15 downto 15) &
  n4(14 downto 14) &
  n4(13 downto 13) &
  n4(12 downto 12) &
  n4(11 downto 11) &
  n4(10 downto 10) &
  n4(9 downto 9) &
  n4(8 downto 8) &
  n4(7 downto 7) &
  n4(6 downto 6) &
  n4(5 downto 5) &
  n4(4 downto 4) &
  n4(3 downto 3) &
  n4(2 downto 2) &
  n4(1 downto 1) &
  n4(0 downto 0);
process (clock_c) begin
  if rising_edge(clock_c) then
    if i5 = "1" then
      n7 <= "0000000000000000";
    elsif i4 = "1" then
      n7 <= n2;
    end if;
  end if;
end process;
process (clock_c) begin
  if rising_edge(clock_c) then
    if i5 = "1" then
      n8 <= "0000000000000000";
    elsif i4 = "1" then
      n8 <= n7;
    end if;
  end if;
end process;
process (clock_c) begin
  if rising_edge(clock_c) then
    if i5 = "1" then
      n9 <= "0000000000000000";
    elsif i4 = "1" then
      n9 <= n3;
    end if;
  end if;
end process;
process (clock_c) begin
  if rising_edge(clock_c) then
    if i5 = "1" then
      n10 <= "0000000000000000";
    elsif i4 = "1" then
      n10 <= n9;
    end if;
  end if;
end process;
process (clock_c) begin
  if rising_edge(clock_c) then 
    if i4 = "1" then
      case i3 is
        when "00" => n11 <= "01111111111111110000000000000000";
        when "01" => n11 <= "01011010100000101010010101111101";
        when "10" => n11 <= "00000000000000001000000000000000";
        when "11" => n11 <= "10100101011111011010010101111101";
        when others => n11 <= "XXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX";
      end case;
    end if;
  end if;
end process;
n12 <= n11(31 downto 31) &
  n11(30 downto 30) &
  n11(29 downto 29) &
  n11(28 downto 28) &
  n11(27 downto 27) &
  n11(26 downto 26) &
  n11(25 downto 25) &
  n11(24 downto 24) &
  n11(23 downto 23) &
  n11(22 downto 22) &
  n11(21 downto 21) &
  n11(20 downto 20) &
  n11(19 downto 19) &
  n11(18 downto 18) &
  n11(17 downto 17) &
  n11(16 downto 16);
n13 <= n11(15 downto 15) &
  n11(14 downto 14) &
  n11(13 downto 13) &
  n11(12 downto 12) &
  n11(11 downto 11) &
  n11(10 downto 10) &
  n11(9 downto 9) &
  n11(8 downto 8) &
  n11(7 downto 7) &
  n11(6 downto 6) &
  n11(5 downto 5) &
  n11(4 downto 4) &
  n11(3 downto 3) &
  n11(2 downto 2) &
  n11(1 downto 1) &
  n11(0 downto 0);
n14 <= unsigned(signed(n5) * signed(n12));
n15 <= n14(30 downto 30) &
  n14(29 downto 29) &
  n14(28 downto 28) &
  n14(27 downto 27) &
  n14(26 downto 26) &
  n14(25 downto 25) &
  n14(24 downto 24) &
  n14(23 downto 23) &
  n14(22 downto 22) &
  n14(21 downto 21) &
  n14(20 downto 20) &
  n14(19 downto 19) &
  n14(18 downto 18) &
  n14(17 downto 17) &
  n14(16 downto 16) &
  n14(15 downto 15);
process (clock_c) begin
  if rising_edge(clock_c) then
    if i5 = "1" then
      n16 <= "0000000000000000";
    elsif i4 = "1" then
      n16 <= n15;
    end if;
  end if;
end process;
n17 <= unsigned(signed(n6) * signed(n13));
n18 <= n17(30 downto 30) &
  n17(29 downto 29) &
  n17(28 downto 28) &
  n17(27 downto 27) &
  n17(26 downto 26) &
  n17(25 downto 25) &
  n17(24 downto 24) &
  n17(23 downto 23) &
  n17(22 downto 22) &
  n17(21 downto 21) &
  n17(20 downto 20) &
  n17(19 downto 19) &
  n17(18 downto 18) &
  n17(17 downto 17) &
  n17(16 downto 16) &
  n17(15 downto 15);
process (clock_c) begin
  if rising_edge(clock_c) then
    if i5 = "1" then
      n19 <= "0000000000000000";
    elsif i4 = "1" then
      n19 <= n18;
    end if;
  end if;
end process;
n20 <= n16 - n19;
process (clock_c) begin
  if rising_edge(clock_c) then
    if i5 = "1" then
      n21 <= "0000000000000000";
    elsif i4 = "1" then
      n21 <= n20;
    end if;
  end if;
end process;
n22 <= unsigned(signed(n5) * signed(n13));
n23 <= n22(30 downto 30) &
  n22(29 downto 29) &
  n22(28 downto 28) &
  n22(27 downto 27) &
  n22(26 downto 26) &
  n22(25 downto 25) &
  n22(24 downto 24) &
  n22(23 downto 23) &
  n22(22 downto 22) &
  n22(21 downto 21) &
  n22(20 downto 20) &
  n22(19 downto 19) &
  n22(18 downto 18) &
  n22(17 downto 17) &
  n22(16 downto 16) &
  n22(15 downto 15);
process (clock_c) begin
  if rising_edge(clock_c) then
    if i5 = "1" then
      n24 <= "0000000000000000";
    elsif i4 = "1" then
      n24 <= n23;
    end if;
  end if;
end process;
n25 <= unsigned(signed(n6) * signed(n12));
n26 <= n25(30 downto 30) &
  n25(29 downto 29) &
  n25(28 downto 28) &
  n25(27 downto 27) &
  n25(26 downto 26) &
  n25(25 downto 25) &
  n25(24 downto 24) &
  n25(23 downto 23) &
  n25(22 downto 22) &
  n25(21 downto 21) &
  n25(20 downto 20) &
  n25(19 downto 19) &
  n25(18 downto 18) &
  n25(17 downto 17) &
  n25(16 downto 16) &
  n25(15 downto 15);
process (clock_c) begin
  if rising_edge(clock_c) then
    if i5 = "1" then
      n27 <= "0000000000000000";
    elsif i4 = "1" then
      n27 <= n26;
    end if;
  end if;
end process;
n28 <= n24 + n27;
process (clock_c) begin
  if rising_edge(clock_c) then
    if i5 = "1" then
      n29 <= "0000000000000000";
    elsif i4 = "1" then
      n29 <= n28;
    end if;
  end if;
end process;
n30 <= n8 + n21;
n31 <= n10 + n29;
n32 <= n30 & n31;
process (clock_c) begin
  if rising_edge(clock_c) then
    if i5 = "1" then
      n33 <= "00000000000000000000000000000000";
    elsif i4 = "1" then
      n33 <= n32;
    end if;
  end if;
end process;
n34 <= n8 - n21;
n35 <= n10 - n29;
n36 <= n34 & n35;
process (clock_c) begin
  if rising_edge(clock_c) then
    if i5 = "1" then
      n37 <= "00000000000000000000000000000000";
    elsif i4 = "1" then
      n37 <= n36;
    end if;
  end if;
end process;
o2 <= n37;
o1 <= n33;
end architecture rtl;

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
entity cf_fft_2048_16_40 is
port (
i1 : in  unsigned(0 downto 0);
i2 : in  unsigned(0 downto 0);
i3 : in  unsigned(0 downto 0);
i4 : in  unsigned(0 downto 0);
i5 : in  unsigned(2 downto 0);
o1 : out unsigned(0 downto 0));
end entity cf_fft_2048_16_40;
architecture rtl of cf_fft_2048_16_40 is
signal n1 : unsigned(2 downto 0);
signal n2 : unsigned(2 downto 0);
signal n3 : unsigned(2 downto 0);
signal n4 : unsigned(0 downto 0);
signal n5 : unsigned(0 downto 0);
signal n6 : unsigned(0 downto 0);
signal n7 : unsigned(0 downto 0);
signal n8 : unsigned(0 downto 0);
signal n9 : unsigned(0 downto 0);
begin
n1 <= "001";
n2 <= "011";
n3 <= "101";
n4 <= "1" when i5 = n1 else "0";
n5 <= "1" when i5 = n2 else "0";
n6 <= "1" when i5 = n3 else "0";
n7 <= i2 when n6 = "1" else i1;
n8 <= i3 when n5 = "1" else n7;
n9 <= i4 when n4 = "1" else n8;
o1 <= n9;
end architecture rtl;

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
entity cf_fft_2048_16_39 is
port (
i1 : in  unsigned(0 downto 0);
i2 : in  unsigned(0 downto 0);
i3 : in  unsigned(0 downto 0);
i4 : in  unsigned(0 downto 0);
i5 : in  unsigned(0 downto 0);
i6 : in  unsigned(0 downto 0);
i7 : in  unsigned(0 downto 0);
i8 : in  unsigned(2 downto 0);
o1 : out unsigned(0 downto 0));
end entity cf_fft_2048_16_39;
architecture rtl of cf_fft_2048_16_39 is
signal n1 : unsigned(2 downto 0);
signal n2 : unsigned(2 downto 0);
signal n3 : unsigned(2 downto 0);
signal n4 : unsigned(0 downto 0);
signal n5 : unsigned(0 downto 0);
signal n6 : unsigned(0 downto 0);
signal n7 : unsigned(0 downto 0);
signal n8 : unsigned(0 downto 0);
signal n9 : unsigned(0 downto 0);
signal s10_1 : unsigned(0 downto 0);
component cf_fft_2048_16_40 is
port (
i1 : in  unsigned(0 downto 0);
i2 : in  unsigned(0 downto 0);
i3 : in  unsigned(0 downto 0);
i4 : in  unsigned(0 downto 0);
i5 : in  unsigned(2 downto 0);
o1 : out unsigned(0 downto 0));
end component cf_fft_2048_16_40;
begin
n1 <= "010";
n2 <= "100";
n3 <= "110";
n4 <= "1" when i8 = n1 else "0";
n5 <= "1" when i8 = n2 else "0";
n6 <= "1" when i8 = n3 else "0";
n7 <= i5 when n6 = "1" else s10_1;
n8 <= i6 when n5 = "1" else n7;
n9 <= i7 when n4 = "1" else n8;
s10 : cf_fft_2048_16_40 port map (i1, i2, i3, i4, i8, s10_1);
o1 <= n9;
end architecture rtl;

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
entity cf_fft_2048_16_38 is
port (
o1 : out unsigned(0 downto 0);
o2 : out unsigned(0 downto 0);
o3 : out unsigned(0 downto 0);
o4 : out unsigned(0 downto 0);
o5 : out unsigned(0 downto 0);
o6 : out unsigned(0 downto 0);
o7 : out unsigned(0 downto 0);
o8 : out unsigned(0 downto 0));
end entity cf_fft_2048_16_38;
architecture rtl of cf_fft_2048_16_38 is
signal n1 : unsigned(0 downto 0);
signal n2 : unsigned(0 downto 0);
signal n3 : unsigned(0 downto 0);
signal n4 : unsigned(0 downto 0);
signal n5 : unsigned(0 downto 0);
signal n6 : unsigned(0 downto 0);
signal n7 : unsigned(0 downto 0);
signal n8 : unsigned(0 downto 0);
begin
n1 <= "0";
n2 <= "1";
n3 <= "0";
n4 <= "1";
n5 <= "0";
n6 <= "1";
n7 <= "0";
n8 <= "0";
o8 <= n8;
o7 <= n7;
o6 <= n6;
o5 <= n5;
o4 <= n4;
o3 <= n3;
o2 <= n2;
o1 <= n1;
end architecture rtl;

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
entity cf_fft_2048_16_37 is
port (
i1 : in  unsigned(0 downto 0);
i2 : in  unsigned(0 downto 0);
i3 : in  unsigned(0 downto 0);
i4 : in  unsigned(2 downto 0);
o1 : out unsigned(0 downto 0));
end entity cf_fft_2048_16_37;
architecture rtl of cf_fft_2048_16_37 is
signal n1 : unsigned(2 downto 0);
signal n2 : unsigned(2 downto 0);
signal n3 : unsigned(2 downto 0);
signal n4 : unsigned(0 downto 0);
signal n5 : unsigned(0 downto 0);
signal n6 : unsigned(0 downto 0);
signal n7 : unsigned(0 downto 0);
signal n8 : unsigned(0 downto 0);
signal n9 : unsigned(0 downto 0);
signal n10 : unsigned(0 downto 0);
begin
n1 <= "010";
n2 <= "100";
n3 <= "110";
n4 <= "1" when i4 = n1 else "0";
n5 <= "1" when i4 = n2 else "0";
n6 <= "1" when i4 = n3 else "0";
n7 <= i1 when n6 = "1" else n10;
n8 <= i2 when n5 = "1" else n7;
n9 <= i3 when n4 = "1" else n8;
n10 <= "1";
o1 <= n9;
end architecture rtl;

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
entity cf_fft_2048_16_36 is
port (
i1 : in  unsigned(2 downto 0);
o1 : out unsigned(0 downto 0));
end entity cf_fft_2048_16_36;
architecture rtl of cf_fft_2048_16_36 is
signal n1 : unsigned(0 downto 0);
signal n2 : unsigned(0 downto 0);
signal n3 : unsigned(0 downto 0);
signal n4 : unsigned(0 downto 0);
signal n5 : unsigned(2 downto 0);
signal n6 : unsigned(0 downto 0);
signal n7 : unsigned(0 downto 0);
signal s8_1 : unsigned(0 downto 0);
component cf_fft_2048_16_37 is
port (
i1 : in  unsigned(0 downto 0);
i2 : in  unsigned(0 downto 0);
i3 : in  unsigned(0 downto 0);
i4 : in  unsigned(2 downto 0);
o1 : out unsigned(0 downto 0));
end component cf_fft_2048_16_37;
begin
n1 <= "0";
n2 <= "0";
n3 <= "0";
n4 <= "0";
n5 <= "000";
n6 <= "1" when i1 = n5 else "0";
n7 <= n4 when n6 = "1" else s8_1;
s8 : cf_fft_2048_16_37 port map (n1, n2, n3, i1, s8_1);
o1 <= n7;
end architecture rtl;

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
entity cf_fft_2048_16_35 is
port (
clock_c : in std_logic;
i1 : in  unsigned(1 downto 0);
i2 : in  unsigned(0 downto 0);
i3 : in  unsigned(0 downto 0);
o1 : out unsigned(0 downto 0));
end entity cf_fft_2048_16_35;
architecture rtl of cf_fft_2048_16_35 is
signal n1 : unsigned(2 downto 0);
signal n2 : unsigned(2 downto 0);
signal n3 : unsigned(0 downto 0);
signal n4 : unsigned(0 downto 0);
signal n5 : unsigned(0 downto 0) := "0";
signal s6_1 : unsigned(0 downto 0);
signal s7_1 : unsigned(0 downto 0);
signal s7_2 : unsigned(0 downto 0);
signal s7_3 : unsigned(0 downto 0);
signal s7_4 : unsigned(0 downto 0);
signal s7_5 : unsigned(0 downto 0);
signal s7_6 : unsigned(0 downto 0);
signal s7_7 : unsigned(0 downto 0);
signal s7_8 : unsigned(0 downto 0);
signal s8_1 : unsigned(0 downto 0);
component cf_fft_2048_16_39 is
port (
i1 : in  unsigned(0 downto 0);
i2 : in  unsigned(0 downto 0);
i3 : in  unsigned(0 downto 0);
i4 : in  unsigned(0 downto 0);
i5 : in  unsigned(0 downto 0);
i6 : in  unsigned(0 downto 0);
i7 : in  unsigned(0 downto 0);
i8 : in  unsigned(2 downto 0);
o1 : out unsigned(0 downto 0));
end component cf_fft_2048_16_39;
component cf_fft_2048_16_38 is
port (
o1 : out unsigned(0 downto 0);
o2 : out unsigned(0 downto 0);
o3 : out unsigned(0 downto 0);
o4 : out unsigned(0 downto 0);
o5 : out unsigned(0 downto 0);
o6 : out unsigned(0 downto 0);
o7 : out unsigned(0 downto 0);
o8 : out unsigned(0 downto 0));
end component cf_fft_2048_16_38;
component cf_fft_2048_16_36 is
port (
i1 : in  unsigned(2 downto 0);
o1 : out unsigned(0 downto 0));
end component cf_fft_2048_16_36;
begin
n1 <= "000";
n2 <= i1 & n5;
n3 <= "1" when n2 = n1 else "0";
n4 <= s7_8 when n3 = "1" else s6_1;
process (clock_c) begin
  if rising_edge(clock_c) then
    if i3 = "1" then
      n5 <= "0";
    elsif i2 = "1" then
      n5 <= n4;
    end if;
  end if;
end process;
s6 : cf_fft_2048_16_39 port map (s7_1, s7_2, s7_3, s7_4, s7_5, s7_6, s7_7, n2, s6_1);
s7 : cf_fft_2048_16_38 port map (s7_1, s7_2, s7_3, s7_4, s7_5, s7_6, s7_7, s7_8);
s8 : cf_fft_2048_16_36 port map (n2, s8_1);
o1 <= s8_1;
end architecture rtl;

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
entity cf_fft_2048_16_34 is
port (
i1 : in  unsigned(0 downto 0);
i2 : in  unsigned(0 downto 0);
i3 : in  unsigned(0 downto 0);
i4 : in  unsigned(0 downto 0);
i5 : in  unsigned(1 downto 0);
o1 : out unsigned(0 downto 0));
end entity cf_fft_2048_16_34;
architecture rtl of cf_fft_2048_16_34 is
signal n1 : unsigned(1 downto 0);
signal n2 : unsigned(1 downto 0);
signal n3 : unsigned(1 downto 0);
signal n4 : unsigned(0 downto 0);
signal n5 : unsigned(0 downto 0);
signal n6 : unsigned(0 downto 0);
signal n7 : unsigned(0 downto 0);
signal n8 : unsigned(0 downto 0);
signal n9 : unsigned(0 downto 0);
begin
n1 <= "00";
n2 <= "10";
n3 <= "01";
n4 <= "1" when i5 = n1 else "0";
n5 <= "1" when i5 = n2 else "0";
n6 <= "1" when i5 = n3 else "0";
n7 <= i2 when n6 = "1" else i1;
n8 <= i3 when n5 = "1" else n7;
n9 <= i4 when n4 = "1" else n8;
o1 <= n9;
end architecture rtl;

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
entity cf_fft_2048_16_33 is
port (
i1 : in  unsigned(1 downto 0);
o1 : out unsigned(0 downto 0));
end entity cf_fft_2048_16_33;
architecture rtl of cf_fft_2048_16_33 is
signal n1 : unsigned(0 downto 0);
signal n2 : unsigned(0 downto 0);
signal n3 : unsigned(1 downto 0);
signal n4 : unsigned(1 downto 0);
signal n5 : unsigned(0 downto 0);
signal n6 : unsigned(0 downto 0);
signal n7 : unsigned(0 downto 0);
signal n8 : unsigned(0 downto 0);
signal n9 : unsigned(0 downto 0);
begin
n1 <= "0";
n2 <= "0";
n3 <= "00";
n4 <= "10";
n5 <= "1" when i1 = n3 else "0";
n6 <= "1" when i1 = n4 else "0";
n7 <= n1 when n6 = "1" else n9;
n8 <= n2 when n5 = "1" else n7;
n9 <= "1";
o1 <= n8;
end architecture rtl;

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
entity cf_fft_2048_16_32 is
port (
clock_c : in std_logic;
i1 : in  unsigned(0 downto 0);
i2 : in  unsigned(0 downto 0);
i3 : in  unsigned(0 downto 0);
o1 : out unsigned(0 downto 0));
end entity cf_fft_2048_16_32;
architecture rtl of cf_fft_2048_16_32 is
signal n1 : unsigned(0 downto 0);
signal n2 : unsigned(0 downto 0);
signal n3 : unsigned(0 downto 0);
signal n4 : unsigned(0 downto 0);
signal n5 : unsigned(1 downto 0);
signal n6 : unsigned(0 downto 0) := "0";
signal s7_1 : unsigned(0 downto 0);
signal s8_1 : unsigned(0 downto 0);
component cf_fft_2048_16_34 is
port (
i1 : in  unsigned(0 downto 0);
i2 : in  unsigned(0 downto 0);
i3 : in  unsigned(0 downto 0);
i4 : in  unsigned(0 downto 0);
i5 : in  unsigned(1 downto 0);
o1 : out unsigned(0 downto 0));
end component cf_fft_2048_16_34;
component cf_fft_2048_16_33 is
port (
i1 : in  unsigned(1 downto 0);
o1 : out unsigned(0 downto 0));
end component cf_fft_2048_16_33;
begin
n1 <= "0";
n2 <= "1";
n3 <= "1";
n4 <= "0";
n5 <= i1 & n6;
process (clock_c) begin
  if rising_edge(clock_c) then
    if i3 = "1" then
      n6 <= "0";
    elsif i2 = "1" then
      n6 <= s7_1;
    end if;
  end if;
end process;
s7 : cf_fft_2048_16_34 port map (n1, n2, n3, n4, n5, s7_1);
s8 : cf_fft_2048_16_33 port map (n5, s8_1);
o1 <= s8_1;
end architecture rtl;

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
entity cf_fft_2048_16_31 is
port (
clock_c : in std_logic;
i1 : in  unsigned(63 downto 0);
i2 : in  unsigned(0 downto 0);
i3 : in  unsigned(8 downto 0);
i4 : in  unsigned(0 downto 0);
i5 : in  unsigned(0 downto 0);
i6 : in  unsigned(0 downto 0);
o1 : out unsigned(63 downto 0));
end entity cf_fft_2048_16_31;
architecture rtl of cf_fft_2048_16_31 is
signal n1 : unsigned(8 downto 0);
signal n2 : unsigned(8 downto 0);
signal n3 : unsigned(8 downto 0) := "000000000";
signal n4 : unsigned(0 downto 0);
signal n5 : unsigned(0 downto 0);
signal n6 : unsigned(63 downto 0);
signal n6a : unsigned(8 downto 0) := "000000000";
type   n6mt is array (511 downto 0) of unsigned(63 downto 0);
signal n6m : n6mt;
signal n7 : unsigned(0 downto 0);
signal n8 : unsigned(63 downto 0);
signal n8a : unsigned(8 downto 0) := "000000000";
type   n8mt is array (511 downto 0) of unsigned(63 downto 0);
signal n8m : n8mt;
signal n9 : unsigned(0 downto 0) := "0";
signal n10 : unsigned(63 downto 0);
signal n11 : unsigned(0 downto 0);
signal s12_1 : unsigned(0 downto 0);
component cf_fft_2048_16_32 is
port (
clock_c : in std_logic;
i1 : in  unsigned(0 downto 0);
i2 : in  unsigned(0 downto 0);
i3 : in  unsigned(0 downto 0);
o1 : out unsigned(0 downto 0));
end component cf_fft_2048_16_32;
begin
n1 <= "000000001";
n2 <= n3 + n1;
process (clock_c) begin
  if rising_edge(clock_c) then
    if n11 = "1" then
      n3 <= "000000000";
    elsif i5 = "1" then
      n3 <= n2;
    end if;
  end if;
end process;
n4 <= not s12_1;
n5 <= i4 and n4;
process (clock_c) begin
  if rising_edge(clock_c) then
    if i5 = "1" then
      if n5 = "1" then
        n6m(to_integer(i3)) <= i1;
      end if;
      n6a <= n3;
    end if;
  end if;
end process;
n6 <= n6m(to_integer(n6a));
n7 <= i4 and s12_1;
process (clock_c) begin
  if rising_edge(clock_c) then
    if i5 = "1" then
      if n7 = "1" then
        n8m(to_integer(i3)) <= i1;
      end if;
      n8a <= n3;
    end if;
  end if;
end process;
n8 <= n8m(to_integer(n8a));
process (clock_c) begin
  if rising_edge(clock_c) then
    if i6 = "1" then
      n9 <= "0";
    elsif i5 = "1" then
      n9 <= n4;
    end if;
  end if;
end process;
n10 <= n8 when n9 = "1" else n6;
n11 <= i2 or i6;
s12 : cf_fft_2048_16_32 port map (clock_c, i2, i5, i6, s12_1);
o1 <= n10;
end architecture rtl;

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
entity cf_fft_2048_16_30 is
port (
clock_c : in std_logic;
i1 : in  unsigned(63 downto 0);
i2 : in  unsigned(0 downto 0);
i3 : in  unsigned(8 downto 0);
i4 : in  unsigned(0 downto 0);
i5 : in  unsigned(0 downto 0);
i6 : in  unsigned(0 downto 0);
o1 : out unsigned(0 downto 0);
o2 : out unsigned(0 downto 0);
o3 : out unsigned(63 downto 0));
end entity cf_fft_2048_16_30;
architecture rtl of cf_fft_2048_16_30 is
signal n1 : unsigned(8 downto 0);
signal n2 : unsigned(8 downto 0);
signal n3 : unsigned(8 downto 0) := "000000000";
signal n4 : unsigned(0 downto 0);
signal n5 : unsigned(0 downto 0) := "0";
signal n6 : unsigned(8 downto 0);
signal n7 : unsigned(0 downto 0);
signal n8 : unsigned(0 downto 0);
signal n9 : unsigned(63 downto 0);
signal n9a : unsigned(8 downto 0) := "000000000";
type   n9mt is array (511 downto 0) of unsigned(63 downto 0);
signal n9m : n9mt;
signal n10 : unsigned(0 downto 0);
signal n11 : unsigned(63 downto 0);
signal n11a : unsigned(8 downto 0) := "000000000";
type   n11mt is array (511 downto 0) of unsigned(63 downto 0);
signal n11m : n11mt;
signal n12 : unsigned(0 downto 0) := "0";
signal n13 : unsigned(63 downto 0);
signal n14 : unsigned(0 downto 0);
signal s15_1 : unsigned(0 downto 0);
component cf_fft_2048_16_32 is
port (
clock_c : in std_logic;
i1 : in  unsigned(0 downto 0);
i2 : in  unsigned(0 downto 0);
i3 : in  unsigned(0 downto 0);
o1 : out unsigned(0 downto 0));
end component cf_fft_2048_16_32;
begin
n1 <= "000000001";
n2 <= n3 + n1;
process (clock_c) begin
  if rising_edge(clock_c) then
    if n14 = "1" then
      n3 <= "000000000";
    elsif i5 = "1" then
      n3 <= n2;
    end if;
  end if;
end process;
n4 <= not s15_1;
process (clock_c) begin
  if rising_edge(clock_c) then
    if i6 = "1" then
      n5 <= "0";
    elsif i5 = "1" then
      n5 <= i2;
    end if;
  end if;
end process;
n6 <= "000000000";
n7 <= "1" when n3 = n6 else "0";
n8 <= i4 and n4;
process (clock_c) begin
  if rising_edge(clock_c) then
    if i5 = "1" then
      if n8 = "1" then
        n9m(to_integer(i3)) <= i1;
      end if;
      n9a <= n3;
    end if;
  end if;
end process;
n9 <= n9m(to_integer(n9a));
n10 <= i4 and s15_1;
process (clock_c) begin
  if rising_edge(clock_c) then
    if i5 = "1" then
      if n10 = "1" then
        n11m(to_integer(i3)) <= i1;
      end if;
      n11a <= n3;
    end if;
  end if;
end process;
n11 <= n11m(to_integer(n11a));
process (clock_c) begin
  if rising_edge(clock_c) then
    if i6 = "1" then
      n12 <= "0";
    elsif i5 = "1" then
      n12 <= n4;
    end if;
  end if;
end process;
n13 <= n11 when n12 = "1" else n9;
n14 <= i2 or i6;
s15 : cf_fft_2048_16_32 port map (clock_c, i2, i5, i6, s15_1);
o3 <= n13;
o2 <= n7;
o1 <= n5;
end architecture rtl;

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
entity cf_fft_2048_16_29 is
port (
i1 : in  unsigned(0 downto 0);
i2 : in  unsigned(0 downto 0);
i3 : in  unsigned(0 downto 0);
i4 : in  unsigned(2 downto 0);
o1 : out unsigned(0 downto 0));
end entity cf_fft_2048_16_29;
architecture rtl of cf_fft_2048_16_29 is
signal n1 : unsigned(2 downto 0);
signal n2 : unsigned(2 downto 0);
signal n3 : unsigned(2 downto 0);
signal n4 : unsigned(0 downto 0);
signal n5 : unsigned(0 downto 0);
signal n6 : unsigned(0 downto 0);
signal n7 : unsigned(0 downto 0);
signal n8 : unsigned(0 downto 0);
signal n9 : unsigned(0 downto 0);
signal n10 : unsigned(0 downto 0);
begin
n1 <= "110";
n2 <= "001";
n3 <= "011";
n4 <= "1" when i4 = n1 else "0";
n5 <= "1" when i4 = n2 else "0";
n6 <= "1" when i4 = n3 else "0";
n7 <= i1 when n6 = "1" else n10;
n8 <= i2 when n5 = "1" else n7;
n9 <= i3 when n4 = "1" else n8;
n10 <= "1";
o1 <= n9;
end architecture rtl;

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
entity cf_fft_2048_16_28 is
port (
i1 : in  unsigned(0 downto 0);
i2 : in  unsigned(0 downto 0);
i3 : in  unsigned(0 downto 0);
i4 : in  unsigned(0 downto 0);
i5 : in  unsigned(0 downto 0);
i6 : in  unsigned(0 downto 0);
i7 : in  unsigned(2 downto 0);
o1 : out unsigned(0 downto 0));
end entity cf_fft_2048_16_28;
architecture rtl of cf_fft_2048_16_28 is
signal n1 : unsigned(2 downto 0);
signal n2 : unsigned(2 downto 0);
signal n3 : unsigned(2 downto 0);
signal n4 : unsigned(0 downto 0);
signal n5 : unsigned(0 downto 0);
signal n6 : unsigned(0 downto 0);
signal n7 : unsigned(0 downto 0);
signal n8 : unsigned(0 downto 0);
signal n9 : unsigned(0 downto 0);
signal s10_1 : unsigned(0 downto 0);
component cf_fft_2048_16_29 is
port (
i1 : in  unsigned(0 downto 0);
i2 : in  unsigned(0 downto 0);
i3 : in  unsigned(0 downto 0);
i4 : in  unsigned(2 downto 0);
o1 : out unsigned(0 downto 0));
end component cf_fft_2048_16_29;
begin
n1 <= "000";
n2 <= "010";
n3 <= "100";
n4 <= "1" when i7 = n1 else "0";
n5 <= "1" when i7 = n2 else "0";
n6 <= "1" when i7 = n3 else "0";
n7 <= i4 when n6 = "1" else s10_1;
n8 <= i5 when n5 = "1" else n7;
n9 <= i6 when n4 = "1" else n8;
s10 : cf_fft_2048_16_29 port map (i1, i2, i3, i7, s10_1);
o1 <= n9;
end architecture rtl;

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
entity cf_fft_2048_16_27 is
port (
clock_c : in std_logic;
i1 : in  unsigned(1 downto 0);
i2 : in  unsigned(0 downto 0);
i3 : in  unsigned(0 downto 0);
o1 : out unsigned(0 downto 0));
end entity cf_fft_2048_16_27;
architecture rtl of cf_fft_2048_16_27 is
signal n1 : unsigned(0 downto 0);
signal n2 : unsigned(0 downto 0);
signal n3 : unsigned(0 downto 0);
signal n4 : unsigned(0 downto 0);
signal n5 : unsigned(0 downto 0);
signal n6 : unsigned(0 downto 0);
signal n7 : unsigned(0 downto 0);
signal n8 : unsigned(0 downto 0);
signal n9 : unsigned(0 downto 0);
signal n10 : unsigned(0 downto 0);
signal n11 : unsigned(0 downto 0);
signal n12 : unsigned(0 downto 0);
signal n13 : unsigned(2 downto 0);
signal n14 : unsigned(0 downto 0) := "0";
signal s15_1 : unsigned(0 downto 0);
signal s16_1 : unsigned(0 downto 0);
component cf_fft_2048_16_28 is
port (
i1 : in  unsigned(0 downto 0);
i2 : in  unsigned(0 downto 0);
i3 : in  unsigned(0 downto 0);
i4 : in  unsigned(0 downto 0);
i5 : in  unsigned(0 downto 0);
i6 : in  unsigned(0 downto 0);
i7 : in  unsigned(2 downto 0);
o1 : out unsigned(0 downto 0));
end component cf_fft_2048_16_28;
begin
n1 <= "0";
n2 <= "1";
n3 <= "1";
n4 <= "1";
n5 <= "0";
n6 <= "0";
n7 <= "0";
n8 <= "1";
n9 <= "1";
n10 <= "1";
n11 <= "0";
n12 <= "0";
n13 <= i1 & n14;
process (clock_c) begin
  if rising_edge(clock_c) then
    if i3 = "1" then
      n14 <= "0";
    elsif i2 = "1" then
      n14 <= s15_1;
    end if;
  end if;
end process;
s15 : cf_fft_2048_16_28 port map (n1, n2, n3, n4, n5, n6, n13, s15_1);
s16 : cf_fft_2048_16_28 port map (n7, n8, n9, n10, n11, n12, n13, s16_1);
o1 <= s16_1;
end architecture rtl;

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
entity cf_fft_2048_16_26 is
port (
clock_c : in std_logic;
i1 : in  unsigned(0 downto 0);
i2 : in  unsigned(0 downto 0);
i3 : in  unsigned(0 downto 0);
o1 : out unsigned(9 downto 0);
o2 : out unsigned(0 downto 0));
end entity cf_fft_2048_16_26;
architecture rtl of cf_fft_2048_16_26 is
signal n1 : unsigned(9 downto 0);
signal n2 : unsigned(9 downto 0);
signal n3 : unsigned(9 downto 0) := "0000000000";
signal n4 : unsigned(9 downto 0);
signal n5 : unsigned(0 downto 0);
signal n6 : unsigned(1 downto 0);
signal n7 : unsigned(0 downto 0) := "0";
signal n8 : unsigned(0 downto 0);
signal n9 : unsigned(0 downto 0);
signal n10 : unsigned(0 downto 0);
signal s11_1 : unsigned(0 downto 0);
component cf_fft_2048_16_27 is
port (
clock_c : in std_logic;
i1 : in  unsigned(1 downto 0);
i2 : in  unsigned(0 downto 0);
i3 : in  unsigned(0 downto 0);
o1 : out unsigned(0 downto 0));
end component cf_fft_2048_16_27;
begin
n1 <= "0000000001";
n2 <= n3 + n1;
process (clock_c) begin
  if rising_edge(clock_c) then
    if n9 = "1" then
      n3 <= "0000000000";
    elsif n10 = "1" then
      n3 <= n2;
    end if;
  end if;
end process;
n4 <= "1111111111";
n5 <= "1" when n3 = n4 else "0";
n6 <= i1 & n5;
process (clock_c) begin
  if rising_edge(clock_c) then
    if i3 = "1" then
      n7 <= "0";
    elsif i2 = "1" then
      n7 <= s11_1;
    end if;
  end if;
end process;
n8 <= n7 and n5;
n9 <= i1 or i3;
n10 <= s11_1 and i2;
s11 : cf_fft_2048_16_27 port map (clock_c, n6, i2, i3, s11_1);
o2 <= n8;
o1 <= n3;
end architecture rtl;

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
entity cf_fft_2048_16_25 is
port (
clock_c : in std_logic;
i1 : in  unsigned(0 downto 0);
i2 : in  unsigned(31 downto 0);
i3 : in  unsigned(31 downto 0);
i4 : in  unsigned(0 downto 0);
i5 : in  unsigned(0 downto 0);
o1 : out unsigned(0 downto 0);
o2 : out unsigned(31 downto 0);
o3 : out unsigned(31 downto 0));
end entity cf_fft_2048_16_25;
architecture rtl of cf_fft_2048_16_25 is
signal n1 : unsigned(1 downto 0);
signal n2 : unsigned(63 downto 0);
signal n3 : unsigned(0 downto 0) := "0";
signal n4 : unsigned(0 downto 0) := "0";
signal n5 : unsigned(0 downto 0) := "0";
signal n6 : unsigned(0 downto 0) := "0";
signal n7 : unsigned(8 downto 0);
signal n8 : unsigned(8 downto 0) := "000000000";
signal n9 : unsigned(8 downto 0) := "000000000";
signal n10 : unsigned(8 downto 0) := "000000000";
signal n11 : unsigned(8 downto 0) := "000000000";
signal n12 : unsigned(0 downto 0);
signal n13 : unsigned(0 downto 0) := "0";
signal n14 : unsigned(0 downto 0) := "0";
signal n15 : unsigned(0 downto 0) := "0";
signal n16 : unsigned(0 downto 0) := "0";
signal n17 : unsigned(0 downto 0);
signal n18 : unsigned(1 downto 0);
signal n19 : unsigned(31 downto 0);
signal n20 : unsigned(31 downto 0);
signal n21 : unsigned(31 downto 0);
signal n22 : unsigned(31 downto 0);
signal n23 : unsigned(31 downto 0);
signal n24 : unsigned(31 downto 0);
signal s25_1 : unsigned(31 downto 0);
signal s25_2 : unsigned(31 downto 0);
signal s26_1 : unsigned(0 downto 0);
signal s27_1 : unsigned(63 downto 0);
signal s28_1 : unsigned(0 downto 0);
signal s28_2 : unsigned(0 downto 0);
signal s28_3 : unsigned(63 downto 0);
signal s29_1 : unsigned(9 downto 0);
signal s29_2 : unsigned(0 downto 0);
component cf_fft_2048_16_41 is
port (
clock_c : in std_logic;
i1 : in  unsigned(31 downto 0);
i2 : in  unsigned(31 downto 0);
i3 : in  unsigned(1 downto 0);
i4 : in  unsigned(0 downto 0);
i5 : in  unsigned(0 downto 0);
o1 : out unsigned(31 downto 0);
o2 : out unsigned(31 downto 0));
end component cf_fft_2048_16_41;
component cf_fft_2048_16_35 is
port (
clock_c : in std_logic;
i1 : in  unsigned(1 downto 0);
i2 : in  unsigned(0 downto 0);
i3 : in  unsigned(0 downto 0);
o1 : out unsigned(0 downto 0));
end component cf_fft_2048_16_35;
component cf_fft_2048_16_31 is
port (
clock_c : in std_logic;
i1 : in  unsigned(63 downto 0);
i2 : in  unsigned(0 downto 0);
i3 : in  unsigned(8 downto 0);
i4 : in  unsigned(0 downto 0);
i5 : in  unsigned(0 downto 0);
i6 : in  unsigned(0 downto 0);
o1 : out unsigned(63 downto 0));
end component cf_fft_2048_16_31;
component cf_fft_2048_16_30 is
port (
clock_c : in std_logic;
i1 : in  unsigned(63 downto 0);
i2 : in  unsigned(0 downto 0);
i3 : in  unsigned(8 downto 0);
i4 : in  unsigned(0 downto 0);
i5 : in  unsigned(0 downto 0);
i6 : in  unsigned(0 downto 0);
o1 : out unsigned(0 downto 0);
o2 : out unsigned(0 downto 0);
o3 : out unsigned(63 downto 0));
end component cf_fft_2048_16_30;
component cf_fft_2048_16_26 is
port (
clock_c : in std_logic;
i1 : in  unsigned(0 downto 0);
i2 : in  unsigned(0 downto 0);
i3 : in  unsigned(0 downto 0);
o1 : out unsigned(9 downto 0);
o2 : out unsigned(0 downto 0));
end component cf_fft_2048_16_26;
begin
n1 <= s29_1(9 downto 9) &
  s29_1(8 downto 8);
n2 <= s25_1 & s25_2;
process (clock_c) begin
  if rising_edge(clock_c) then
    if i5 = "1" then
      n3 <= "0";
    elsif i4 = "1" then
      n3 <= s29_2;
    end if;
  end if;
end process;
process (clock_c) begin
  if rising_edge(clock_c) then
    if i5 = "1" then
      n4 <= "0";
    elsif i4 = "1" then
      n4 <= n3;
    end if;
  end if;
end process;
process (clock_c) begin
  if rising_edge(clock_c) then
    if i5 = "1" then
      n5 <= "0";
    elsif i4 = "1" then
      n5 <= n4;
    end if;
  end if;
end process;
process (clock_c) begin
  if rising_edge(clock_c) then
    if i5 = "1" then
      n6 <= "0";
    elsif i4 = "1" then
      n6 <= n5;
    end if;
  end if;
end process;
n7 <= s29_1(9 downto 9) &
  s29_1(8 downto 8) &
  s29_1(7 downto 7) &
  s29_1(6 downto 6) &
  s29_1(5 downto 5) &
  s29_1(4 downto 4) &
  s29_1(3 downto 3) &
  s29_1(2 downto 2) &
  s29_1(1 downto 1);
process (clock_c) begin
  if rising_edge(clock_c) then
    if i5 = "1" then
      n8 <= "000000000";
    elsif i4 = "1" then
      n8 <= n7;
    end if;
  end if;
end process;
process (clock_c) begin
  if rising_edge(clock_c) then
    if i5 = "1" then
      n9 <= "000000000";
    elsif i4 = "1" then
      n9 <= n8;
    end if;
  end if;
end process;
process (clock_c) begin
  if rising_edge(clock_c) then
    if i5 = "1" then
      n10 <= "000000000";
    elsif i4 = "1" then
      n10 <= n9;
    end if;
  end if;
end process;
process (clock_c) begin
  if rising_edge(clock_c) then
    if i5 = "1" then
      n11 <= "000000000";
    elsif i4 = "1" then
      n11 <= n10;
    end if;
  end if;
end process;
n12 <= s29_1(0 downto 0);
process (clock_c) begin
  if rising_edge(clock_c) then
    if i5 = "1" then
      n13 <= "0";
    elsif i4 = "1" then
      n13 <= n12;
    end if;
  end if;
end process;
process (clock_c) begin
  if rising_edge(clock_c) then
    if i5 = "1" then
      n14 <= "0";
    elsif i4 = "1" then
      n14 <= n13;
    end if;
  end if;
end process;
process (clock_c) begin
  if rising_edge(clock_c) then
    if i5 = "1" then
      n15 <= "0";
    elsif i4 = "1" then
      n15 <= n14;
    end if;
  end if;
end process;
process (clock_c) begin
  if rising_edge(clock_c) then
    if i5 = "1" then
      n16 <= "0";
    elsif i4 = "1" then
      n16 <= n15;
    end if;
  end if;
end process;
n17 <= not n16;
n18 <= s28_2 & s28_1;
n19 <= s28_3(63 downto 63) &
  s28_3(62 downto 62) &
  s28_3(61 downto 61) &
  s28_3(60 downto 60) &
  s28_3(59 downto 59) &
  s28_3(58 downto 58) &
  s28_3(57 downto 57) &
  s28_3(56 downto 56) &
  s28_3(55 downto 55) &
  s28_3(54 downto 54) &
  s28_3(53 downto 53) &
  s28_3(52 downto 52) &
  s28_3(51 downto 51) &
  s28_3(50 downto 50) &
  s28_3(49 downto 49) &
  s28_3(48 downto 48) &
  s28_3(47 downto 47) &
  s28_3(46 downto 46) &
  s28_3(45 downto 45) &
  s28_3(44 downto 44) &
  s28_3(43 downto 43) &
  s28_3(42 downto 42) &
  s28_3(41 downto 41) &
  s28_3(40 downto 40) &
  s28_3(39 downto 39) &
  s28_3(38 downto 38) &
  s28_3(37 downto 37) &
  s28_3(36 downto 36) &
  s28_3(35 downto 35) &
  s28_3(34 downto 34) &
  s28_3(33 downto 33) &
  s28_3(32 downto 32);
n20 <= s28_3(31 downto 31) &
  s28_3(30 downto 30) &
  s28_3(29 downto 29) &
  s28_3(28 downto 28) &
  s28_3(27 downto 27) &
  s28_3(26 downto 26) &
  s28_3(25 downto 25) &
  s28_3(24 downto 24) &
  s28_3(23 downto 23) &
  s28_3(22 downto 22) &
  s28_3(21 downto 21) &
  s28_3(20 downto 20) &
  s28_3(19 downto 19) &
  s28_3(18 downto 18) &
  s28_3(17 downto 17) &
  s28_3(16 downto 16) &
  s28_3(15 downto 15) &
  s28_3(14 downto 14) &
  s28_3(13 downto 13) &
  s28_3(12 downto 12) &
  s28_3(11 downto 11) &
  s28_3(10 downto 10) &
  s28_3(9 downto 9) &
  s28_3(8 downto 8) &
  s28_3(7 downto 7) &
  s28_3(6 downto 6) &
  s28_3(5 downto 5) &
  s28_3(4 downto 4) &
  s28_3(3 downto 3) &
  s28_3(2 downto 2) &
  s28_3(1 downto 1) &
  s28_3(0 downto 0);
n21 <= s27_1(63 downto 63) &
  s27_1(62 downto 62) &
  s27_1(61 downto 61) &
  s27_1(60 downto 60) &
  s27_1(59 downto 59) &
  s27_1(58 downto 58) &
  s27_1(57 downto 57) &
  s27_1(56 downto 56) &
  s27_1(55 downto 55) &
  s27_1(54 downto 54) &
  s27_1(53 downto 53) &
  s27_1(52 downto 52) &
  s27_1(51 downto 51) &
  s27_1(50 downto 50) &
  s27_1(49 downto 49) &
  s27_1(48 downto 48) &
  s27_1(47 downto 47) &
  s27_1(46 downto 46) &
  s27_1(45 downto 45) &
  s27_1(44 downto 44) &
  s27_1(43 downto 43) &
  s27_1(42 downto 42) &
  s27_1(41 downto 41) &
  s27_1(40 downto 40) &
  s27_1(39 downto 39) &
  s27_1(38 downto 38) &
  s27_1(37 downto 37) &
  s27_1(36 downto 36) &
  s27_1(35 downto 35) &
  s27_1(34 downto 34) &
  s27_1(33 downto 33) &
  s27_1(32 downto 32);
n22 <= s27_1(31 downto 31) &
  s27_1(30 downto 30) &
  s27_1(29 downto 29) &
  s27_1(28 downto 28) &
  s27_1(27 downto 27) &
  s27_1(26 downto 26) &
  s27_1(25 downto 25) &
  s27_1(24 downto 24) &
  s27_1(23 downto 23) &
  s27_1(22 downto 22) &
  s27_1(21 downto 21) &
  s27_1(20 downto 20) &
  s27_1(19 downto 19) &
  s27_1(18 downto 18) &
  s27_1(17 downto 17) &
  s27_1(16 downto 16) &
  s27_1(15 downto 15) &
  s27_1(14 downto 14) &
  s27_1(13 downto 13) &
  s27_1(12 downto 12) &
  s27_1(11 downto 11) &
  s27_1(10 downto 10) &
  s27_1(9 downto 9) &
  s27_1(8 downto 8) &
  s27_1(7 downto 7) &
  s27_1(6 downto 6) &
  s27_1(5 downto 5) &
  s27_1(4 downto 4) &
  s27_1(3 downto 3) &
  s27_1(2 downto 2) &
  s27_1(1 downto 1) &
  s27_1(0 downto 0);
n23 <= n20 when s26_1 = "1" else n19;
n24 <= n22 when s26_1 = "1" else n21;
s25 : cf_fft_2048_16_41 port map (clock_c, i2, i3, n1, i4, i5, s25_1, s25_2);
s26 : cf_fft_2048_16_35 port map (clock_c, n18, i4, i5, s26_1);
s27 : cf_fft_2048_16_31 port map (clock_c, n2, n6, n11, n16, i4, i5, s27_1);
s28 : cf_fft_2048_16_30 port map (clock_c, n2, n6, n11, n17, i4, i5, s28_1, s28_2, s28_3);
s29 : cf_fft_2048_16_26 port map (clock_c, i1, i4, i5, s29_1, s29_2);
o3 <= n24;
o2 <= n23;
o1 <= s28_1;
end architecture rtl;

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
entity cf_fft_2048_16_24 is
port (
clock_c : in std_logic;
i1 : in  unsigned(31 downto 0);
i2 : in  unsigned(31 downto 0);
i3 : in  unsigned(9 downto 0);
i4 : in  unsigned(0 downto 0);
i5 : in  unsigned(0 downto 0);
o1 : out unsigned(31 downto 0);
o2 : out unsigned(31 downto 0));
end entity cf_fft_2048_16_24;
architecture rtl of cf_fft_2048_16_24 is
signal n1 : unsigned(31 downto 0) := "00000000000000000000000000000000";
signal n2 : unsigned(15 downto 0);
signal n3 : unsigned(15 downto 0);
signal n4 : unsigned(31 downto 0) := "00000000000000000000000000000000";
signal n5 : unsigned(15 downto 0);
signal n6 : unsigned(15 downto 0);
signal n7 : unsigned(15 downto 0) := "0000000000000000";
signal n8 : unsigned(15 downto 0) := "0000000000000000";
signal n9 : unsigned(15 downto 0) := "0000000000000000";
signal n10 : unsigned(15 downto 0) := "0000000000000000";
signal n11 : unsigned(31 downto 0) := "00000000000000000000000000000000";
signal n12 : unsigned(15 downto 0);
signal n13 : unsigned(15 downto 0);
signal n14 : unsigned(31 downto 0);
signal n15 : unsigned(15 downto 0);
signal n16 : unsigned(15 downto 0) := "0000000000000000";
signal n17 : unsigned(31 downto 0);
signal n18 : unsigned(15 downto 0);
signal n19 : unsigned(15 downto 0) := "0000000000000000";
signal n20 : unsigned(15 downto 0);
signal n21 : unsigned(15 downto 0) := "0000000000000000";
signal n22 : unsigned(31 downto 0);
signal n23 : unsigned(15 downto 0);
signal n24 : unsigned(15 downto 0) := "0000000000000000";
signal n25 : unsigned(31 downto 0);
signal n26 : unsigned(15 downto 0);
signal n27 : unsigned(15 downto 0) := "0000000000000000";
signal n28 : unsigned(15 downto 0);
signal n29 : unsigned(15 downto 0) := "0000000000000000";
signal n30 : unsigned(15 downto 0);
signal n31 : unsigned(15 downto 0);
signal n32 : unsigned(31 downto 0);
signal n33 : unsigned(31 downto 0) := "00000000000000000000000000000000";
signal n34 : unsigned(15 downto 0);
signal n35 : unsigned(15 downto 0);
signal n36 : unsigned(31 downto 0);
signal n37 : unsigned(31 downto 0) := "00000000000000000000000000000000";
begin
process (clock_c) begin
  if rising_edge(clock_c) then
    if i5 = "1" then
      n1 <= "00000000000000000000000000000000";
    elsif i4 = "1" then
      n1 <= i1;
    end if;
  end if;
end process;
n2 <= n1(31 downto 31) &
  n1(30 downto 30) &
  n1(29 downto 29) &
  n1(28 downto 28) &
  n1(27 downto 27) &
  n1(26 downto 26) &
  n1(25 downto 25) &
  n1(24 downto 24) &
  n1(23 downto 23) &
  n1(22 downto 22) &
  n1(21 downto 21) &
  n1(20 downto 20) &
  n1(19 downto 19) &
  n1(18 downto 18) &
  n1(17 downto 17) &
  n1(16 downto 16);
n3 <= n1(15 downto 15) &
  n1(14 downto 14) &
  n1(13 downto 13) &
  n1(12 downto 12) &
  n1(11 downto 11) &
  n1(10 downto 10) &
  n1(9 downto 9) &
  n1(8 downto 8) &
  n1(7 downto 7) &
  n1(6 downto 6) &
  n1(5 downto 5) &
  n1(4 downto 4) &
  n1(3 downto 3) &
  n1(2 downto 2) &
  n1(1 downto 1) &
  n1(0 downto 0);
process (clock_c) begin
  if rising_edge(clock_c) then
    if i5 = "1" then
      n4 <= "00000000000000000000000000000000";
    elsif i4 = "1" then
      n4 <= i2;
    end if;
  end if;
end process;
n5 <= n4(31 downto 31) &
  n4(30 downto 30) &
  n4(29 downto 29) &
  n4(28 downto 28) &
  n4(27 downto 27) &
  n4(26 downto 26) &
  n4(25 downto 25) &
  n4(24 downto 24) &
  n4(23 downto 23) &
  n4(22 downto 22) &
  n4(21 downto 21) &
  n4(20 downto 20) &
  n4(19 downto 19) &
  n4(18 downto 18) &
  n4(17 downto 17) &
  n4(16 downto 16);
n6 <= n4(15 downto 15) &
  n4(14 downto 14) &
  n4(13 downto 13) &
  n4(12 downto 12) &
  n4(11 downto 11) &
  n4(10 downto 10) &
  n4(9 downto 9) &
  n4(8 downto 8) &
  n4(7 downto 7) &
  n4(6 downto 6) &
  n4(5 downto 5) &
  n4(4 downto 4) &
  n4(3 downto 3) &
  n4(2 downto 2) &
  n4(1 downto 1) &
  n4(0 downto 0);
process (clock_c) begin
  if rising_edge(clock_c) then
    if i5 = "1" then
      n7 <= "0000000000000000";
    elsif i4 = "1" then
      n7 <= n2;
    end if;
  end if;
end process;
process (clock_c) begin
  if rising_edge(clock_c) then
    if i5 = "1" then
      n8 <= "0000000000000000";
    elsif i4 = "1" then
      n8 <= n7;
    end if;
  end if;
end process;
process (clock_c) begin
  if rising_edge(clock_c) then
    if i5 = "1" then
      n9 <= "0000000000000000";
    elsif i4 = "1" then
      n9 <= n3;
    end if;
  end if;
end process;
process (clock_c) begin
  if rising_edge(clock_c) then
    if i5 = "1" then
      n10 <= "0000000000000000";
    elsif i4 = "1" then
      n10 <= n9;
    end if;
  end if;
end process;
process (clock_c) begin
  if rising_edge(clock_c) then 
    if i4 = "1" then
      case i3 is
        when "0000000000" => n11 <= "01111111111111110000000000000000";
        when "0000000001" => n11 <= "01111111111111111111111110011011";
        when "0000000010" => n11 <= "01111111111111111111111100110110";
        when "0000000011" => n11 <= "01111111111111101111111011010010";
        when "0000000100" => n11 <= "01111111111111011111111001101101";
        when "0000000101" => n11 <= "01111111111111001111111000001001";
        when "0000000110" => n11 <= "01111111111110101111110110100100";
        when "0000000111" => n11 <= "01111111111110001111110101000000";
        when "0000001000" => n11 <= "01111111111101101111110011011011";
        when "0000001001" => n11 <= "01111111111100111111110001110111";
        when "0000001010" => n11 <= "01111111111100001111110000010010";
        when "0000001011" => n11 <= "01111111111011011111101110101110";
        when "0000001100" => n11 <= "01111111111010011111101101001001";
        when "0000001101" => n11 <= "01111111111001011111101011100101";
        when "0000001110" => n11 <= "01111111111000011111101010000000";
        when "0000001111" => n11 <= "01111111110111011111101000011100";
        when "0000010000" => n11 <= "01111111110110001111100110111000";
        when "0000010001" => n11 <= "01111111110100111111100101010011";
        when "0000010010" => n11 <= "01111111110011101111100011101111";
        when "0000010011" => n11 <= "01111111110010001111100010001010";
        when "0000010100" => n11 <= "01111111110000101111100000100110";
        when "0000010101" => n11 <= "01111111101111001111011111000010";
        when "0000010110" => n11 <= "01111111101101011111011101011101";
        when "0000010111" => n11 <= "01111111101011101111011011111001";
        when "0000011000" => n11 <= "01111111101001111111011010010101";
        when "0000011001" => n11 <= "01111111100111111111011000110001";
        when "0000011010" => n11 <= "01111111100101111111010111001100";
        when "0000011011" => n11 <= "01111111100011111111010101101000";
        when "0000011100" => n11 <= "01111111100001111111010100000100";
        when "0000011101" => n11 <= "01111111011111101111010010100000";
        when "0000011110" => n11 <= "01111111011101011111010000111100";
        when "0000011111" => n11 <= "01111111011010111111001111011000";
        when "0000100000" => n11 <= "01111111011000101111001101110100";
        when "0000100001" => n11 <= "01111111010110001111001100010000";
        when "0000100010" => n11 <= "01111111010011011111001010101100";
        when "0000100011" => n11 <= "01111111010000111111001001001000";
        when "0000100100" => n11 <= "01111111001110001111000111100100";
        when "0000100101" => n11 <= "01111111001011011111000110000000";
        when "0000100110" => n11 <= "01111111001000011111000100011100";
        when "0000100111" => n11 <= "01111111000101011111000010111000";
        when "0000101000" => n11 <= "01111111000010011111000001010100";
        when "0000101001" => n11 <= "01111110111111011110111111110001";
        when "0000101010" => n11 <= "01111110111100001110111110001101";
        when "0000101011" => n11 <= "01111110111000111110111100101001";
        when "0000101100" => n11 <= "01111110110101011110111011000110";
        when "0000101101" => n11 <= "01111110110010001110111001100010";
        when "0000101110" => n11 <= "01111110101110101110110111111110";
        when "0000101111" => n11 <= "01111110101010111110110110011011";
        when "0000110000" => n11 <= "01111110100111011110110100110111";
        when "0000110001" => n11 <= "01111110100011101110110011010100";
        when "0000110010" => n11 <= "01111110011111111110110001110001";
        when "0000110011" => n11 <= "01111110011011111110110000001101";
        when "0000110100" => n11 <= "01111110010111111110101110101010";
        when "0000110101" => n11 <= "01111110010011111110101101000111";
        when "0000110110" => n11 <= "01111110001111111110101011100100";
        when "0000110111" => n11 <= "01111110001011101110101010000000";
        when "0000111000" => n11 <= "01111110000111011110101000011101";
        when "0000111001" => n11 <= "01111110000011001110100110111010";
        when "0000111010" => n11 <= "01111101111110101110100101010111";
        when "0000111011" => n11 <= "01111101111010001110100011110101";
        when "0000111100" => n11 <= "01111101110101101110100010010010";
        when "0000111101" => n11 <= "01111101110000111110100000101111";
        when "0000111110" => n11 <= "01111101101100001110011111001100";
        when "0000111111" => n11 <= "01111101100111011110011101101001";
        when "0001000000" => n11 <= "01111101100010101110011100000111";
        when "0001000001" => n11 <= "01111101011101101110011010100100";
        when "0001000010" => n11 <= "01111101011000101110011001000010";
        when "0001000011" => n11 <= "01111101010011101110010111011111";
        when "0001000100" => n11 <= "01111101001110011110010101111101";
        when "0001000101" => n11 <= "01111101001001001110010100011011";
        when "0001000110" => n11 <= "01111101000011111110010010111000";
        when "0001000111" => n11 <= "01111100111110011110010001010110";
        when "0001001000" => n11 <= "01111100111000111110001111110100";
        when "0001001001" => n11 <= "01111100110011011110001110010010";
        when "0001001010" => n11 <= "01111100101101111110001100110000";
        when "0001001011" => n11 <= "01111100101000001110001011001110";
        when "0001001100" => n11 <= "01111100100010011110001001101100";
        when "0001001101" => n11 <= "01111100011100011110001000001010";
        when "0001001110" => n11 <= "01111100010110101110000110101001";
        when "0001001111" => n11 <= "01111100010000101110000101000111";
        when "0001010000" => n11 <= "01111100001010011110000011100110";
        when "0001010001" => n11 <= "01111100000100011110000010000100";
        when "0001010010" => n11 <= "01111011111110001110000000100011";
        when "0001010011" => n11 <= "01111011110111111101111111000001";
        when "0001010100" => n11 <= "01111011110001011101111101100000";
        when "0001010101" => n11 <= "01111011101011001101111011111111";
        when "0001010110" => n11 <= "01111011100100101101111010011110";
        when "0001010111" => n11 <= "01111011011101111101111000111101";
        when "0001011000" => n11 <= "01111011010111011101110111011100";
        when "0001011001" => n11 <= "01111011010000101101110101111011";
        when "0001011010" => n11 <= "01111011001001101101110100011010";
        when "0001011011" => n11 <= "01111011000010111101110010111010";
        when "0001011100" => n11 <= "01111010111011111101110001011001";
        when "0001011101" => n11 <= "01111010110100111101101111111000";
        when "0001011110" => n11 <= "01111010101101101101101110011000";
        when "0001011111" => n11 <= "01111010100110101101101100111000";
        when "0001100000" => n11 <= "01111010011111011101101011010111";
        when "0001100001" => n11 <= "01111010010111111101101001110111";
        when "0001100010" => n11 <= "01111010010000101101101000010111";
        when "0001100011" => n11 <= "01111010001001001101100110110111";
        when "0001100100" => n11 <= "01111010000001011101100101010111";
        when "0001100101" => n11 <= "01111001111001111101100011111000";
        when "0001100110" => n11 <= "01111001110010001101100010011000";
        when "0001100111" => n11 <= "01111001101010011101100000111000";
        when "0001101000" => n11 <= "01111001100010101101011111011001";
        when "0001101001" => n11 <= "01111001011010101101011101111001";
        when "0001101010" => n11 <= "01111001010010101101011100011010";
        when "0001101011" => n11 <= "01111001001010101101011010111011";
        when "0001101100" => n11 <= "01111001000010011101011001011100";
        when "0001101101" => n11 <= "01111000111010001101010111111101";
        when "0001101110" => n11 <= "01111000110001111101010110011110";
        when "0001101111" => n11 <= "01111000101001101101010100111111";
        when "0001110000" => n11 <= "01111000100001001101010011100000";
        when "0001110001" => n11 <= "01111000011000101101010010000010";
        when "0001110010" => n11 <= "01111000010000001101010000100011";
        when "0001110011" => n11 <= "01111000000111011101001111000101";
        when "0001110100" => n11 <= "01110111111110101101001101100111";
        when "0001110101" => n11 <= "01110111110101111101001100001000";
        when "0001110110" => n11 <= "01110111101101001101001010101010";
        when "0001110111" => n11 <= "01110111100100001101001001001100";
        when "0001111000" => n11 <= "01110111011011001101000111101110";
        when "0001111001" => n11 <= "01110111010001111101000110010001";
        when "0001111010" => n11 <= "01110111001000111101000100110011";
        when "0001111011" => n11 <= "01110110111111101101000011010110";
        when "0001111100" => n11 <= "01110110110110011101000001111000";
        when "0001111101" => n11 <= "01110110101100111101000000011011";
        when "0001111110" => n11 <= "01110110100011101100111110111110";
        when "0001111111" => n11 <= "01110110011010001100111101100001";
        when "0010000000" => n11 <= "01110110010000011100111100000100";
        when "0010000001" => n11 <= "01110110000110111100111010100111";
        when "0010000010" => n11 <= "01110101111101001100111001001010";
        when "0010000011" => n11 <= "01110101110011001100110111101110";
        when "0010000100" => n11 <= "01110101101001011100110110010001";
        when "0010000101" => n11 <= "01110101011111011100110100110101";
        when "0010000110" => n11 <= "01110101010101011100110011011001";
        when "0010000111" => n11 <= "01110101001011011100110001111101";
        when "0010001000" => n11 <= "01110101000001001100110000100001";
        when "0010001001" => n11 <= "01110100110110111100101111000101";
        when "0010001010" => n11 <= "01110100101100101100101101101001";
        when "0010001011" => n11 <= "01110100100010011100101100001101";
        when "0010001100" => n11 <= "01110100010111111100101010110010";
        when "0010001101" => n11 <= "01110100001101011100101001010111";
        when "0010001110" => n11 <= "01110100000010111100100111111011";
        when "0010001111" => n11 <= "01110011111000001100100110100000";
        when "0010010000" => n11 <= "01110011101101011100100101000101";
        when "0010010001" => n11 <= "01110011100010101100100011101011";
        when "0010010010" => n11 <= "01110011010111111100100010010000";
        when "0010010011" => n11 <= "01110011001100111100100000110101";
        when "0010010100" => n11 <= "01110011000001111100011111011011";
        when "0010010101" => n11 <= "01110010110110111100011110000001";
        when "0010010110" => n11 <= "01110010101011111100011100100111";
        when "0010010111" => n11 <= "01110010100000101100011011001101";
        when "0010011000" => n11 <= "01110010010101011100011001110011";
        when "0010011001" => n11 <= "01110010001001111100011000011001";
        when "0010011010" => n11 <= "01110001111110101100010110111111";
        when "0010011011" => n11 <= "01110001110011001100010101100110";
        when "0010011100" => n11 <= "01110001100111101100010100001101";
        when "0010011101" => n11 <= "01110001011011111100010010110011";
        when "0010011110" => n11 <= "01110001010000011100010001011010";
        when "0010011111" => n11 <= "01110001000100101100010000000010";
        when "0010100000" => n11 <= "01110000111000101100001110101001";
        when "0010100001" => n11 <= "01110000101100111100001101010000";
        when "0010100010" => n11 <= "01110000100000111100001011111000";
        when "0010100011" => n11 <= "01110000010100111100001010011111";
        when "0010100100" => n11 <= "01110000001000111100001001000111";
        when "0010100101" => n11 <= "01101111111100101100000111101111";
        when "0010100110" => n11 <= "01101111110000011100000110010111";
        when "0010100111" => n11 <= "01101111100100001100000101000000";
        when "0010101000" => n11 <= "01101111010111111100000011101000";
        when "0010101001" => n11 <= "01101111001011011100000010010001";
        when "0010101010" => n11 <= "01101110111110111100000000111010";
        when "0010101011" => n11 <= "01101110110010011011111111100010";
        when "0010101100" => n11 <= "01101110100101101011111110001100";
        when "0010101101" => n11 <= "01101110011000111011111100110101";
        when "0010101110" => n11 <= "01101110001100001011111011011110";
        when "0010101111" => n11 <= "01101101111111011011111010001000";
        when "0010110000" => n11 <= "01101101110010101011111000110001";
        when "0010110001" => n11 <= "01101101100101101011110111011011";
        when "0010110010" => n11 <= "01101101011000101011110110000101";
        when "0010110011" => n11 <= "01101101001011011011110100101111";
        when "0010110100" => n11 <= "01101100111110011011110011011010";
        when "0010110101" => n11 <= "01101100110001001011110010000100";
        when "0010110110" => n11 <= "01101100100011111011110000101111";
        when "0010110111" => n11 <= "01101100010110011011101111011010";
        when "0010111000" => n11 <= "01101100001001001011101110000101";
        when "0010111001" => n11 <= "01101011111011101011101100110000";
        when "0010111010" => n11 <= "01101011101110001011101011011011";
        when "0010111011" => n11 <= "01101011100000011011101010000111";
        when "0010111100" => n11 <= "01101011010010101011101000110010";
        when "0010111101" => n11 <= "01101011000100111011100111011110";
        when "0010111110" => n11 <= "01101010110111001011100110001010";
        when "0010111111" => n11 <= "01101010101001011011100100110110";
        when "0011000000" => n11 <= "01101010011011011011100011100011";
        when "0011000001" => n11 <= "01101010001101011011100010001111";
        when "0011000010" => n11 <= "01101001111111011011100000111100";
        when "0011000011" => n11 <= "01101001110001001011011111101001";
        when "0011000100" => n11 <= "01101001100011001011011110010110";
        when "0011000101" => n11 <= "01101001010100111011011101000011";
        when "0011000110" => n11 <= "01101001000110011011011011110000";
        when "0011000111" => n11 <= "01101000111000001011011010011110";
        when "0011001000" => n11 <= "01101000101001101011011001001011";
        when "0011001001" => n11 <= "01101000011011001011010111111001";
        when "0011001010" => n11 <= "01101000001100101011010110100111";
        when "0011001011" => n11 <= "01100111111101111011010101010110";
        when "0011001100" => n11 <= "01100111101111011011010100000100";
        when "0011001101" => n11 <= "01100111100000101011010010110011";
        when "0011001110" => n11 <= "01100111010001101011010001100001";
        when "0011001111" => n11 <= "01100111000010111011010000010000";
        when "0011010000" => n11 <= "01100110110011111011001111000000";
        when "0011010001" => n11 <= "01100110100100111011001101101111";
        when "0011010010" => n11 <= "01100110010101111011001100011110";
        when "0011010011" => n11 <= "01100110000110101011001011001110";
        when "0011010100" => n11 <= "01100101110111011011001001111110";
        when "0011010101" => n11 <= "01100101101000001011001000101110";
        when "0011010110" => n11 <= "01100101011000111011000111011110";
        when "0011010111" => n11 <= "01100101001001101011000110001111";
        when "0011011000" => n11 <= "01100100111010001011000101000000";
        when "0011011001" => n11 <= "01100100101010101011000011110000";
        when "0011011010" => n11 <= "01100100011011001011000010100001";
        when "0011011011" => n11 <= "01100100001011011011000001010011";
        when "0011011100" => n11 <= "01100011111011111011000000000100";
        when "0011011101" => n11 <= "01100011101100001010111110110110";
        when "0011011110" => n11 <= "01100011011100011010111101101000";
        when "0011011111" => n11 <= "01100011001100011010111100011010";
        when "0011100000" => n11 <= "01100010111100101010111011001100";
        when "0011100001" => n11 <= "01100010101100101010111001111110";
        when "0011100010" => n11 <= "01100010011100011010111000110001";
        when "0011100011" => n11 <= "01100010001100011010110111100011";
        when "0011100100" => n11 <= "01100001111100011010110110010110";
        when "0011100101" => n11 <= "01100001101100001010110101001010";
        when "0011100110" => n11 <= "01100001011011111010110011111101";
        when "0011100111" => n11 <= "01100001001011011010110010110001";
        when "0011101000" => n11 <= "01100000111011001010110001100100";
        when "0011101001" => n11 <= "01100000101010101010110000011000";
        when "0011101010" => n11 <= "01100000011010001010101111001100";
        when "0011101011" => n11 <= "01100000001001101010101110000001";
        when "0011101100" => n11 <= "01011111111000111010101100110101";
        when "0011101101" => n11 <= "01011111101000001010101011101010";
        when "0011101110" => n11 <= "01011111010111101010101010011111";
        when "0011101111" => n11 <= "01011111000110101010101001010100";
        when "0011110000" => n11 <= "01011110110101111010101000001010";
        when "0011110001" => n11 <= "01011110100100111010100110111111";
        when "0011110010" => n11 <= "01011110010100001010100101110101";
        when "0011110011" => n11 <= "01011110000010111010100100101011";
        when "0011110100" => n11 <= "01011101110001111010100011100010";
        when "0011110101" => n11 <= "01011101100000111010100010011000";
        when "0011110110" => n11 <= "01011101001111101010100001001111";
        when "0011110111" => n11 <= "01011100111110011010100000000110";
        when "0011111000" => n11 <= "01011100101101001010011110111101";
        when "0011111001" => n11 <= "01011100011011101010011101110100";
        when "0011111010" => n11 <= "01011100001010011010011100101011";
        when "0011111011" => n11 <= "01011011111000111010011011100011";
        when "0011111100" => n11 <= "01011011100111011010011010011011";
        when "0011111101" => n11 <= "01011011010101101010011001010011";
        when "0011111110" => n11 <= "01011011000100001010011000001100";
        when "0011111111" => n11 <= "01011010110010011010010111000100";
        when "0100000000" => n11 <= "01011010100000101010010101111101";
        when "0100000001" => n11 <= "01011010001110111010010100110110";
        when "0100000010" => n11 <= "01011001111100111010010011101111";
        when "0100000011" => n11 <= "01011001101011001010010010101001";
        when "0100000100" => n11 <= "01011001011001001010010001100010";
        when "0100000101" => n11 <= "01011001000111001010010000011100";
        when "0100000110" => n11 <= "01011000110101001010001111010110";
        when "0100000111" => n11 <= "01011000100010111010001110010001";
        when "0100001000" => n11 <= "01011000010000101010001101001011";
        when "0100001001" => n11 <= "01010111111110011010001100000110";
        when "0100001010" => n11 <= "01010111101100001010001011000001";
        when "0100001011" => n11 <= "01010111011001111010001001111100";
        when "0100001100" => n11 <= "01010111000111011010001000111000";
        when "0100001101" => n11 <= "01010110110101001010000111110100";
        when "0100001110" => n11 <= "01010110100010101010000110101111";
        when "0100001111" => n11 <= "01010110010000001010000101101100";
        when "0100010000" => n11 <= "01010101111101011010000100101000";
        when "0100010001" => n11 <= "01010101101010111010000011100101";
        when "0100010010" => n11 <= "01010101011000001010000010100001";
        when "0100010011" => n11 <= "01010101000101011010000001011111";
        when "0100010100" => n11 <= "01010100110010101010000000011100";
        when "0100010101" => n11 <= "01010100011111101001111111011001";
        when "0100010110" => n11 <= "01010100001100111001111110010111";
        when "0100010111" => n11 <= "01010011111001111001111101010101";
        when "0100011000" => n11 <= "01010011100110111001111100010011";
        when "0100011001" => n11 <= "01010011010011101001111011010010";
        when "0100011010" => n11 <= "01010011000000101001111010010000";
        when "0100011011" => n11 <= "01010010101101011001111001001111";
        when "0100011100" => n11 <= "01010010011010011001111000001110";
        when "0100011101" => n11 <= "01010010000111001001110111001110";
        when "0100011110" => n11 <= "01010001110011101001110110001110";
        when "0100011111" => n11 <= "01010001100000011001110101001101";
        when "0100100000" => n11 <= "01010001001100111001110100001101";
        when "0100100001" => n11 <= "01010000111001011001110011001110";
        when "0100100010" => n11 <= "01010000100101111001110010001110";
        when "0100100011" => n11 <= "01010000010010011001110001001111";
        when "0100100100" => n11 <= "01001111111110111001110000010000";
        when "0100100101" => n11 <= "01001111101011001001101111010010";
        when "0100100110" => n11 <= "01001111010111101001101110010011";
        when "0100100111" => n11 <= "01001111000011111001101101010101";
        when "0100101000" => n11 <= "01001110101111111001101100010111";
        when "0100101001" => n11 <= "01001110011100001001101011011001";
        when "0100101010" => n11 <= "01001110001000011001101010011100";
        when "0100101011" => n11 <= "01001101110100011001101001011111";
        when "0100101100" => n11 <= "01001101100000011001101000100010";
        when "0100101101" => n11 <= "01001101001100011001100111100101";
        when "0100101110" => n11 <= "01001100111000011001100110101000";
        when "0100101111" => n11 <= "01001100100100001001100101101100";
        when "0100110000" => n11 <= "01001100001111111001100100110000";
        when "0100110001" => n11 <= "01001011111011111001100011110100";
        when "0100110010" => n11 <= "01001011100111101001100010111001";
        when "0100110011" => n11 <= "01001011010011001001100001111101";
        when "0100110100" => n11 <= "01001010111110111001100001000010";
        when "0100110101" => n11 <= "01001010101010011001100000001000";
        when "0100110110" => n11 <= "01001010010110001001011111001101";
        when "0100110111" => n11 <= "01001010000001101001011110010011";
        when "0100111000" => n11 <= "01001001101101001001011101011001";
        when "0100111001" => n11 <= "01001001011000011001011100011111";
        when "0100111010" => n11 <= "01001001000011111001011011100110";
        when "0100111011" => n11 <= "01001000101111001001011010101100";
        when "0100111100" => n11 <= "01001000011010011001011001110011";
        when "0100111101" => n11 <= "01001000000101101001011000111011";
        when "0100111110" => n11 <= "01000111110000111001011000000010";
        when "0100111111" => n11 <= "01000111011100001001010111001010";
        when "0101000000" => n11 <= "01000111000111001001010110010010";
        when "0101000001" => n11 <= "01000110110010011001010101011010";
        when "0101000010" => n11 <= "01000110011101011001010100100011";
        when "0101000011" => n11 <= "01000110001000011001010011101100";
        when "0101000100" => n11 <= "01000101110011011001010010110101";
        when "0101000101" => n11 <= "01000101011110001001010001111110";
        when "0101000110" => n11 <= "01000101001001001001010001000111";
        when "0101000111" => n11 <= "01000100110011111001010000010001";
        when "0101001000" => n11 <= "01000100011110101001001111011011";
        when "0101001001" => n11 <= "01000100001001011001001110100110";
        when "0101001010" => n11 <= "01000011110100001001001101110000";
        when "0101001011" => n11 <= "01000011011110111001001100111011";
        when "0101001100" => n11 <= "01000011001001011001001100000110";
        when "0101001101" => n11 <= "01000010110100001001001011010010";
        when "0101001110" => n11 <= "01000010011110101001001010011101";
        when "0101001111" => n11 <= "01000010001001001001001001101001";
        when "0101010000" => n11 <= "01000001110011101001001000110101";
        when "0101010001" => n11 <= "01000001011101111001001000000010";
        when "0101010010" => n11 <= "01000001001000011001000111001111";
        when "0101010011" => n11 <= "01000000110010101001000110011100";
        when "0101010100" => n11 <= "01000000011100111001000101101001";
        when "0101010101" => n11 <= "01000000000111011001000100110110";
        when "0101010110" => n11 <= "00111111110001011001000100000100";
        when "0101010111" => n11 <= "00111111011011101001000011010010";
        when "0101011000" => n11 <= "00111111000101111001000010100000";
        when "0101011001" => n11 <= "00111110101111111001000001101111";
        when "0101011010" => n11 <= "00111110011010001001000000111110";
        when "0101011011" => n11 <= "00111110000100001001000000001101";
        when "0101011100" => n11 <= "00111101101110001000111111011100";
        when "0101011101" => n11 <= "00111101011000001000111110101100";
        when "0101011110" => n11 <= "00111101000001111000111101111100";
        when "0101011111" => n11 <= "00111100101011111000111101001100";
        when "0101100000" => n11 <= "00111100010101101000111100011101";
        when "0101100001" => n11 <= "00111011111111011000111011101101";
        when "0101100010" => n11 <= "00111011101001011000111010111110";
        when "0101100011" => n11 <= "00111011010011001000111010010000";
        when "0101100100" => n11 <= "00111010111100101000111001100001";
        when "0101100101" => n11 <= "00111010100110011000111000110011";
        when "0101100110" => n11 <= "00111010010000001000111000000101";
        when "0101100111" => n11 <= "00111001111001101000110111011000";
        when "0101101000" => n11 <= "00111001100011001000110110101010";
        when "0101101001" => n11 <= "00111001001100101000110101111101";
        when "0101101010" => n11 <= "00111000110110001000110101010000";
        when "0101101011" => n11 <= "00111000011111101000110100100100";
        when "0101101100" => n11 <= "00111000001001001000110011111000";
        when "0101101101" => n11 <= "00110111110010101000110011001100";
        when "0101101110" => n11 <= "00110111011011111000110010100000";
        when "0101101111" => n11 <= "00110111000101001000110001110101";
        when "0101110000" => n11 <= "00110110101110101000110001001010";
        when "0101110001" => n11 <= "00110110010111111000110000011111";
        when "0101110010" => n11 <= "00110110000001001000101111110100";
        when "0101110011" => n11 <= "00110101101010001000101111001010";
        when "0101110100" => n11 <= "00110101010011011000101110100000";
        when "0101110101" => n11 <= "00110100111100101000101101110110";
        when "0101110110" => n11 <= "00110100100101101000101101001101";
        when "0101110111" => n11 <= "00110100001110101000101100100100";
        when "0101111000" => n11 <= "00110011110111101000101011111011";
        when "0101111001" => n11 <= "00110011100000101000101011010010";
        when "0101111010" => n11 <= "00110011001001101000101010101010";
        when "0101111011" => n11 <= "00110010110010101000101010000010";
        when "0101111100" => n11 <= "00110010011011101000101001011010";
        when "0101111101" => n11 <= "00110010000100011000101000110011";
        when "0101111110" => n11 <= "00110001101101011000101000001011";
        when "0101111111" => n11 <= "00110001010110001000100111100100";
        when "0110000000" => n11 <= "00110000111110111000100110111110";
        when "0110000001" => n11 <= "00110000100111101000100110010111";
        when "0110000010" => n11 <= "00110000010000011000100101110001";
        when "0110000011" => n11 <= "00101111111001001000100101001100";
        when "0110000100" => n11 <= "00101111100001111000100100100110";
        when "0110000101" => n11 <= "00101111001010011000100100000001";
        when "0110000110" => n11 <= "00101110110011001000100011011100";
        when "0110000111" => n11 <= "00101110011011101000100010111000";
        when "0110001000" => n11 <= "00101110000100011000100010010011";
        when "0110001001" => n11 <= "00101101101100111000100001101111";
        when "0110001010" => n11 <= "00101101010101011000100001001011";
        when "0110001011" => n11 <= "00101100111101111000100000101000";
        when "0110001100" => n11 <= "00101100100110001000100000000101";
        when "0110001101" => n11 <= "00101100001110101000011111100010";
        when "0110001110" => n11 <= "00101011110111001000011110111111";
        when "0110001111" => n11 <= "00101011011111011000011110011101";
        when "0110010000" => n11 <= "00101011000111111000011101111011";
        when "0110010001" => n11 <= "00101010110000001000011101011001";
        when "0110010010" => n11 <= "00101010011000011000011100111000";
        when "0110010011" => n11 <= "00101010000000101000011100010111";
        when "0110010100" => n11 <= "00101001101000111000011011110110";
        when "0110010101" => n11 <= "00101001010001001000011011010101";
        when "0110010110" => n11 <= "00101000111001011000011010110101";
        when "0110010111" => n11 <= "00101000100001101000011010010101";
        when "0110011000" => n11 <= "00101000001001101000011001110101";
        when "0110011001" => n11 <= "00100111110001111000011001010110";
        when "0110011010" => n11 <= "00100111011001111000011000110111";
        when "0110011011" => n11 <= "00100111000001111000011000011000";
        when "0110011100" => n11 <= "00100110101010001000010111111010";
        when "0110011101" => n11 <= "00100110010010001000010111011011";
        when "0110011110" => n11 <= "00100101111010001000010110111101";
        when "0110011111" => n11 <= "00100101100010001000010110100000";
        when "0110100000" => n11 <= "00100101001010001000010110000010";
        when "0110100001" => n11 <= "00100100110001111000010101100101";
        when "0110100010" => n11 <= "00100100011001111000010101001001";
        when "0110100011" => n11 <= "00100100000001111000010100101100";
        when "0110100100" => n11 <= "00100011101001101000010100010000";
        when "0110100101" => n11 <= "00100011010001011000010011110100";
        when "0110100110" => n11 <= "00100010111001011000010011011001";
        when "0110100111" => n11 <= "00100010100001001000010010111101";
        when "0110101000" => n11 <= "00100010001000111000010010100010";
        when "0110101001" => n11 <= "00100001110000101000010010001000";
        when "0110101010" => n11 <= "00100001011000011000010001101101";
        when "0110101011" => n11 <= "00100001000000001000010001010011";
        when "0110101100" => n11 <= "00100000100111111000010000111010";
        when "0110101101" => n11 <= "00100000001111101000010000100000";
        when "0110101110" => n11 <= "00011111110111001000010000000111";
        when "0110101111" => n11 <= "00011111011110111000001111101110";
        when "0110110000" => n11 <= "00011111000110011000001111010110";
        when "0110110001" => n11 <= "00011110101110001000001110111101";
        when "0110110010" => n11 <= "00011110010101101000001110100101";
        when "0110110011" => n11 <= "00011101111101011000001110001110";
        when "0110110100" => n11 <= "00011101100100111000001101110110";
        when "0110110101" => n11 <= "00011101001100011000001101011111";
        when "0110110110" => n11 <= "00011100110011111000001101001000";
        when "0110110111" => n11 <= "00011100011011011000001100110010";
        when "0110111000" => n11 <= "00011100000010111000001100011100";
        when "0110111001" => n11 <= "00011011101010011000001100000110";
        when "0110111010" => n11 <= "00011011010001111000001011110000";
        when "0110111011" => n11 <= "00011010111001001000001011011011";
        when "0110111100" => n11 <= "00011010100000101000001011000110";
        when "0110111101" => n11 <= "00011010001000001000001010110001";
        when "0110111110" => n11 <= "00011001101111011000001010011101";
        when "0110111111" => n11 <= "00011001010110111000001010001001";
        when "0111000000" => n11 <= "00011000111110001000001001110101";
        when "0111000001" => n11 <= "00011000100101101000001001100010";
        when "0111000010" => n11 <= "00011000001100111000001001001111";
        when "0111000011" => n11 <= "00010111110100001000001000111100";
        when "0111000100" => n11 <= "00010111011011011000001000101001";
        when "0111000101" => n11 <= "00010111000010101000001000010111";
        when "0111000110" => n11 <= "00010110101010001000001000000101";
        when "0111000111" => n11 <= "00010110010001011000000111110011";
        when "0111001000" => n11 <= "00010101111000101000000111100010";
        when "0111001001" => n11 <= "00010101011111111000000111010001";
        when "0111001010" => n11 <= "00010101000110111000000111000000";
        when "0111001011" => n11 <= "00010100101110001000000110110000";
        when "0111001100" => n11 <= "00010100010101011000000110100000";
        when "0111001101" => n11 <= "00010011111100101000000110010000";
        when "0111001110" => n11 <= "00010011100011101000000110000000";
        when "0111001111" => n11 <= "00010011001010111000000101110001";
        when "0111010000" => n11 <= "00010010110010001000000101100010";
        when "0111010001" => n11 <= "00010010011001001000000101010100";
        when "0111010010" => n11 <= "00010010000000011000000101000101";
        when "0111010011" => n11 <= "00010001100111011000000100110111";
        when "0111010100" => n11 <= "00010001001110011000000100101010";
        when "0111010101" => n11 <= "00010000110101101000000100011100";
        when "0111010110" => n11 <= "00010000011100101000000100001111";
        when "0111010111" => n11 <= "00010000000011101000000100000010";
        when "0111011000" => n11 <= "00001111101010111000000011110110";
        when "0111011001" => n11 <= "00001111010001111000000011101010";
        when "0111011010" => n11 <= "00001110111000111000000011011110";
        when "0111011011" => n11 <= "00001110011111111000000011010010";
        when "0111011100" => n11 <= "00001110000110111000000011000111";
        when "0111011101" => n11 <= "00001101101101111000000010111100";
        when "0111011110" => n11 <= "00001101010100111000000010110010";
        when "0111011111" => n11 <= "00001100111011111000000010100111";
        when "0111100000" => n11 <= "00001100100010111000000010011101";
        when "0111100001" => n11 <= "00001100001001111000000010010100";
        when "0111100010" => n11 <= "00001011110000111000000010001010";
        when "0111100011" => n11 <= "00001011010111111000000010000001";
        when "0111100100" => n11 <= "00001010111110111000000001111000";
        when "0111100101" => n11 <= "00001010100101111000000001110000";
        when "0111100110" => n11 <= "00001010001100111000000001101000";
        when "0111100111" => n11 <= "00001001110011101000000001100000";
        when "0111101000" => n11 <= "00001001011010101000000001011000";
        when "0111101001" => n11 <= "00001001000001101000000001010001";
        when "0111101010" => n11 <= "00001000101000101000000001001010";
        when "0111101011" => n11 <= "00001000001111011000000001000011";
        when "0111101100" => n11 <= "00000111110110011000000000111101";
        when "0111101101" => n11 <= "00000111011101011000000000110111";
        when "0111101110" => n11 <= "00000111000100001000000000110001";
        when "0111101111" => n11 <= "00000110101011001000000000101100";
        when "0111110000" => n11 <= "00000110010001111000000000100111";
        when "0111110001" => n11 <= "00000101111000111000000000100010";
        when "0111110010" => n11 <= "00000101011111111000000000011110";
        when "0111110011" => n11 <= "00000101000110101000000000011010";
        when "0111110100" => n11 <= "00000100101101101000000000010110";
        when "0111110101" => n11 <= "00000100010100011000000000010010";
        when "0111110110" => n11 <= "00000011111011011000000000001111";
        when "0111110111" => n11 <= "00000011100010001000000000001100";
        when "0111111000" => n11 <= "00000011001001001000000000001001";
        when "0111111001" => n11 <= "00000010101111111000000000000111";
        when "0111111010" => n11 <= "00000010010110111000000000000101";
        when "0111111011" => n11 <= "00000001111101101000000000000011";
        when "0111111100" => n11 <= "00000001100100101000000000000010";
        when "0111111101" => n11 <= "00000001001011011000000000000001";
        when "0111111110" => n11 <= "00000000110010011000000000000000";
        when "0111111111" => n11 <= "00000000011001001000000000000000";
        when "1000000000" => n11 <= "00000000000000001000000000000000";
        when "1000000001" => n11 <= "11111111100110111000000000000000";
        when "1000000010" => n11 <= "11111111001101101000000000000000";
        when "1000000011" => n11 <= "11111110110100101000000000000001";
        when "1000000100" => n11 <= "11111110011011011000000000000010";
        when "1000000101" => n11 <= "11111110000010011000000000000011";
        when "1000000110" => n11 <= "11111101101001001000000000000101";
        when "1000000111" => n11 <= "11111101010000001000000000000111";
        when "1000001000" => n11 <= "11111100110110111000000000001001";
        when "1000001001" => n11 <= "11111100011101111000000000001100";
        when "1000001010" => n11 <= "11111100000100101000000000001111";
        when "1000001011" => n11 <= "11111011101011101000000000010010";
        when "1000001100" => n11 <= "11111011010010011000000000010110";
        when "1000001101" => n11 <= "11111010111001011000000000011010";
        when "1000001110" => n11 <= "11111010100000001000000000011110";
        when "1000001111" => n11 <= "11111010000111001000000000100010";
        when "1000010000" => n11 <= "11111001101110001000000000100111";
        when "1000010001" => n11 <= "11111001010100111000000000101100";
        when "1000010010" => n11 <= "11111000111011111000000000110001";
        when "1000010011" => n11 <= "11111000100010101000000000110111";
        when "1000010100" => n11 <= "11111000001001101000000000111101";
        when "1000010101" => n11 <= "11110111110000101000000001000011";
        when "1000010110" => n11 <= "11110111010111011000000001001010";
        when "1000010111" => n11 <= "11110110111110011000000001010001";
        when "1000011000" => n11 <= "11110110100101011000000001011000";
        when "1000011001" => n11 <= "11110110001100011000000001100000";
        when "1000011010" => n11 <= "11110101110011001000000001101000";
        when "1000011011" => n11 <= "11110101011010001000000001110000";
        when "1000011100" => n11 <= "11110101000001001000000001111000";
        when "1000011101" => n11 <= "11110100101000001000000010000001";
        when "1000011110" => n11 <= "11110100001111001000000010001010";
        when "1000011111" => n11 <= "11110011110110001000000010010100";
        when "1000100000" => n11 <= "11110011011101001000000010011101";
        when "1000100001" => n11 <= "11110011000100001000000010100111";
        when "1000100010" => n11 <= "11110010101011001000000010110010";
        when "1000100011" => n11 <= "11110010010010001000000010111100";
        when "1000100100" => n11 <= "11110001111001001000000011000111";
        when "1000100101" => n11 <= "11110001100000001000000011010010";
        when "1000100110" => n11 <= "11110001000111001000000011011110";
        when "1000100111" => n11 <= "11110000101110001000000011101010";
        when "1000101000" => n11 <= "11110000010101001000000011110110";
        when "1000101001" => n11 <= "11101111111100011000000100000010";
        when "1000101010" => n11 <= "11101111100011011000000100001111";
        when "1000101011" => n11 <= "11101111001010011000000100011100";
        when "1000101100" => n11 <= "11101110110001101000000100101010";
        when "1000101101" => n11 <= "11101110011000101000000100110111";
        when "1000101110" => n11 <= "11101101111111101000000101000101";
        when "1000101111" => n11 <= "11101101100110111000000101010100";
        when "1000110000" => n11 <= "11101101001101111000000101100010";
        when "1000110001" => n11 <= "11101100110101001000000101110001";
        when "1000110010" => n11 <= "11101100011100011000000110000000";
        when "1000110011" => n11 <= "11101100000011011000000110010000";
        when "1000110100" => n11 <= "11101011101010101000000110100000";
        when "1000110101" => n11 <= "11101011010001111000000110110000";
        when "1000110110" => n11 <= "11101010111001001000000111000000";
        when "1000110111" => n11 <= "11101010100000001000000111010001";
        when "1000111000" => n11 <= "11101010000111011000000111100010";
        when "1000111001" => n11 <= "11101001101110101000000111110011";
        when "1000111010" => n11 <= "11101001010101111000001000000101";
        when "1000111011" => n11 <= "11101000111101011000001000010111";
        when "1000111100" => n11 <= "11101000100100101000001000101001";
        when "1000111101" => n11 <= "11101000001011111000001000111100";
        when "1000111110" => n11 <= "11100111110011001000001001001111";
        when "1000111111" => n11 <= "11100111011010011000001001100010";
        when "1001000000" => n11 <= "11100111000001111000001001110101";
        when "1001000001" => n11 <= "11100110101001001000001010001001";
        when "1001000010" => n11 <= "11100110010000101000001010011101";
        when "1001000011" => n11 <= "11100101110111111000001010110001";
        when "1001000100" => n11 <= "11100101011111011000001011000110";
        when "1001000101" => n11 <= "11100101000110111000001011011011";
        when "1001000110" => n11 <= "11100100101110001000001011110000";
        when "1001000111" => n11 <= "11100100010101101000001100000110";
        when "1001001000" => n11 <= "11100011111101001000001100011100";
        when "1001001001" => n11 <= "11100011100100101000001100110010";
        when "1001001010" => n11 <= "11100011001100001000001101001000";
        when "1001001011" => n11 <= "11100010110011101000001101011111";
        when "1001001100" => n11 <= "11100010011011001000001101110110";
        when "1001001101" => n11 <= "11100010000010101000001110001110";
        when "1001001110" => n11 <= "11100001101010011000001110100101";
        when "1001001111" => n11 <= "11100001010001111000001110111101";
        when "1001010000" => n11 <= "11100000111001101000001111010110";
        when "1001010001" => n11 <= "11100000100001001000001111101110";
        when "1001010010" => n11 <= "11100000001000111000010000000111";
        when "1001010011" => n11 <= "11011111110000011000010000100000";
        when "1001010100" => n11 <= "11011111011000001000010000111010";
        when "1001010101" => n11 <= "11011110111111111000010001010011";
        when "1001010110" => n11 <= "11011110100111101000010001101101";
        when "1001010111" => n11 <= "11011110001111011000010010001000";
        when "1001011000" => n11 <= "11011101110111001000010010100010";
        when "1001011001" => n11 <= "11011101011110111000010010111101";
        when "1001011010" => n11 <= "11011101000110101000010011011001";
        when "1001011011" => n11 <= "11011100101110101000010011110100";
        when "1001011100" => n11 <= "11011100010110011000010100010000";
        when "1001011101" => n11 <= "11011011111110001000010100101100";
        when "1001011110" => n11 <= "11011011100110001000010101001001";
        when "1001011111" => n11 <= "11011011001110001000010101100101";
        when "1001100000" => n11 <= "11011010110101111000010110000010";
        when "1001100001" => n11 <= "11011010011101111000010110100000";
        when "1001100010" => n11 <= "11011010000101111000010110111101";
        when "1001100011" => n11 <= "11011001101101111000010111011011";
        when "1001100100" => n11 <= "11011001010101111000010111111010";
        when "1001100101" => n11 <= "11011000111110001000011000011000";
        when "1001100110" => n11 <= "11011000100110001000011000110111";
        when "1001100111" => n11 <= "11011000001110001000011001010110";
        when "1001101000" => n11 <= "11010111110110011000011001110101";
        when "1001101001" => n11 <= "11010111011110011000011010010101";
        when "1001101010" => n11 <= "11010111000110101000011010110101";
        when "1001101011" => n11 <= "11010110101110111000011011010101";
        when "1001101100" => n11 <= "11010110010111001000011011110110";
        when "1001101101" => n11 <= "11010101111111011000011100010111";
        when "1001101110" => n11 <= "11010101100111101000011100111000";
        when "1001101111" => n11 <= "11010101001111111000011101011001";
        when "1001110000" => n11 <= "11010100111000001000011101111011";
        when "1001110001" => n11 <= "11010100100000101000011110011101";
        when "1001110010" => n11 <= "11010100001000111000011110111111";
        when "1001110011" => n11 <= "11010011110001011000011111100010";
        when "1001110100" => n11 <= "11010011011001111000100000000101";
        when "1001110101" => n11 <= "11010011000010001000100000101000";
        when "1001110110" => n11 <= "11010010101010101000100001001011";
        when "1001110111" => n11 <= "11010010010011001000100001101111";
        when "1001111000" => n11 <= "11010001111011101000100010010011";
        when "1001111001" => n11 <= "11010001100100011000100010111000";
        when "1001111010" => n11 <= "11010001001100111000100011011100";
        when "1001111011" => n11 <= "11010000110101101000100100000001";
        when "1001111100" => n11 <= "11010000011110001000100100100110";
        when "1001111101" => n11 <= "11010000000110111000100101001100";
        when "1001111110" => n11 <= "11001111101111101000100101110001";
        when "1001111111" => n11 <= "11001111011000011000100110010111";
        when "1010000000" => n11 <= "11001111000001001000100110111110";
        when "1010000001" => n11 <= "11001110101001111000100111100100";
        when "1010000010" => n11 <= "11001110010010101000101000001011";
        when "1010000011" => n11 <= "11001101111011101000101000110011";
        when "1010000100" => n11 <= "11001101100100011000101001011010";
        when "1010000101" => n11 <= "11001101001101011000101010000010";
        when "1010000110" => n11 <= "11001100110110011000101010101010";
        when "1010000111" => n11 <= "11001100011111011000101011010010";
        when "1010001000" => n11 <= "11001100001000011000101011111011";
        when "1010001001" => n11 <= "11001011110001011000101100100100";
        when "1010001010" => n11 <= "11001011011010011000101101001101";
        when "1010001011" => n11 <= "11001011000011011000101101110110";
        when "1010001100" => n11 <= "11001010101100101000101110100000";
        when "1010001101" => n11 <= "11001010010101111000101111001010";
        when "1010001110" => n11 <= "11001001111110111000101111110100";
        when "1010001111" => n11 <= "11001001101000001000110000011111";
        when "1010010000" => n11 <= "11001001010001011000110001001010";
        when "1010010001" => n11 <= "11001000111010111000110001110101";
        when "1010010010" => n11 <= "11001000100100001000110010100000";
        when "1010010011" => n11 <= "11001000001101011000110011001100";
        when "1010010100" => n11 <= "11000111110110111000110011111000";
        when "1010010101" => n11 <= "11000111100000011000110100100100";
        when "1010010110" => n11 <= "11000111001001111000110101010000";
        when "1010010111" => n11 <= "11000110110011011000110101111101";
        when "1010011000" => n11 <= "11000110011100111000110110101010";
        when "1010011001" => n11 <= "11000110000110011000110111011000";
        when "1010011010" => n11 <= "11000101101111111000111000000101";
        when "1010011011" => n11 <= "11000101011001101000111000110011";
        when "1010011100" => n11 <= "11000101000011011000111001100001";
        when "1010011101" => n11 <= "11000100101100111000111010010000";
        when "1010011110" => n11 <= "11000100010110101000111010111110";
        when "1010011111" => n11 <= "11000100000000101000111011101101";
        when "1010100000" => n11 <= "11000011101010011000111100011101";
        when "1010100001" => n11 <= "11000011010100001000111101001100";
        when "1010100010" => n11 <= "11000010111110001000111101111100";
        when "1010100011" => n11 <= "11000010100111111000111110101100";
        when "1010100100" => n11 <= "11000010010001111000111111011100";
        when "1010100101" => n11 <= "11000001111011111001000000001101";
        when "1010100110" => n11 <= "11000001100101111001000000111110";
        when "1010100111" => n11 <= "11000001010000001001000001101111";
        when "1010101000" => n11 <= "11000000111010001001000010100000";
        when "1010101001" => n11 <= "11000000100100011001000011010010";
        when "1010101010" => n11 <= "11000000001110101001000100000100";
        when "1010101011" => n11 <= "10111111111000101001000100110110";
        when "1010101100" => n11 <= "10111111100011001001000101101001";
        when "1010101101" => n11 <= "10111111001101011001000110011100";
        when "1010101110" => n11 <= "10111110110111101001000111001111";
        when "1010101111" => n11 <= "10111110100010001001001000000010";
        when "1010110000" => n11 <= "10111110001100011001001000110101";
        when "1010110001" => n11 <= "10111101110110111001001001101001";
        when "1010110010" => n11 <= "10111101100001011001001010011101";
        when "1010110011" => n11 <= "10111101001011111001001011010010";
        when "1010110100" => n11 <= "10111100110110101001001100000110";
        when "1010110101" => n11 <= "10111100100001001001001100111011";
        when "1010110110" => n11 <= "10111100001011111001001101110000";
        when "1010110111" => n11 <= "10111011110110101001001110100110";
        when "1010111000" => n11 <= "10111011100001011001001111011011";
        when "1010111001" => n11 <= "10111011001100001001010000010001";
        when "1010111010" => n11 <= "10111010110110111001010001000111";
        when "1010111011" => n11 <= "10111010100001111001010001111110";
        when "1010111100" => n11 <= "10111010001100101001010010110101";
        when "1010111101" => n11 <= "10111001110111101001010011101100";
        when "1010111110" => n11 <= "10111001100010101001010100100011";
        when "1010111111" => n11 <= "10111001001101101001010101011010";
        when "1011000000" => n11 <= "10111000111000111001010110010010";
        when "1011000001" => n11 <= "10111000100011111001010111001010";
        when "1011000010" => n11 <= "10111000001111001001011000000010";
        when "1011000011" => n11 <= "10110111111010011001011000111011";
        when "1011000100" => n11 <= "10110111100101101001011001110011";
        when "1011000101" => n11 <= "10110111010000111001011010101100";
        when "1011000110" => n11 <= "10110110111100001001011011100110";
        when "1011000111" => n11 <= "10110110100111101001011100011111";
        when "1011001000" => n11 <= "10110110010010111001011101011001";
        when "1011001001" => n11 <= "10110101111110011001011110010011";
        when "1011001010" => n11 <= "10110101101001111001011111001101";
        when "1011001011" => n11 <= "10110101010101101001100000001000";
        when "1011001100" => n11 <= "10110101000001001001100001000010";
        when "1011001101" => n11 <= "10110100101100111001100001111101";
        when "1011001110" => n11 <= "10110100011000011001100010111001";
        when "1011001111" => n11 <= "10110100000100001001100011110100";
        when "1011010000" => n11 <= "10110011110000001001100100110000";
        when "1011010001" => n11 <= "10110011011011111001100101101100";
        when "1011010010" => n11 <= "10110011000111101001100110101000";
        when "1011010011" => n11 <= "10110010110011101001100111100101";
        when "1011010100" => n11 <= "10110010011111101001101000100010";
        when "1011010101" => n11 <= "10110010001011101001101001011111";
        when "1011010110" => n11 <= "10110001110111101001101010011100";
        when "1011010111" => n11 <= "10110001100011111001101011011001";
        when "1011011000" => n11 <= "10110001010000001001101100010111";
        when "1011011001" => n11 <= "10110000111100001001101101010101";
        when "1011011010" => n11 <= "10110000101000011001101110010011";
        when "1011011011" => n11 <= "10110000010100111001101111010010";
        when "1011011100" => n11 <= "10110000000001001001110000010000";
        when "1011011101" => n11 <= "10101111101101101001110001001111";
        when "1011011110" => n11 <= "10101111011010001001110010001110";
        when "1011011111" => n11 <= "10101111000110101001110011001110";
        when "1011100000" => n11 <= "10101110110011001001110100001101";
        when "1011100001" => n11 <= "10101110011111101001110101001101";
        when "1011100010" => n11 <= "10101110001100011001110110001110";
        when "1011100011" => n11 <= "10101101111000111001110111001110";
        when "1011100100" => n11 <= "10101101100101101001111000001110";
        when "1011100101" => n11 <= "10101101010010101001111001001111";
        when "1011100110" => n11 <= "10101100111111011001111010010000";
        when "1011100111" => n11 <= "10101100101100011001111011010010";
        when "1011101000" => n11 <= "10101100011001001001111100010011";
        when "1011101001" => n11 <= "10101100000110001001111101010101";
        when "1011101010" => n11 <= "10101011110011001001111110010111";
        when "1011101011" => n11 <= "10101011100000011001111111011001";
        when "1011101100" => n11 <= "10101011001101011010000000011100";
        when "1011101101" => n11 <= "10101010111010101010000001011111";
        when "1011101110" => n11 <= "10101010100111111010000010100001";
        when "1011101111" => n11 <= "10101010010101001010000011100101";
        when "1011110000" => n11 <= "10101010000010101010000100101000";
        when "1011110001" => n11 <= "10101001101111111010000101101100";
        when "1011110010" => n11 <= "10101001011101011010000110101111";
        when "1011110011" => n11 <= "10101001001010111010000111110100";
        when "1011110100" => n11 <= "10101000111000101010001000111000";
        when "1011110101" => n11 <= "10101000100110001010001001111100";
        when "1011110110" => n11 <= "10101000010011111010001011000001";
        when "1011110111" => n11 <= "10101000000001101010001100000110";
        when "1011111000" => n11 <= "10100111101111011010001101001011";
        when "1011111001" => n11 <= "10100111011101001010001110010001";
        when "1011111010" => n11 <= "10100111001010111010001111010110";
        when "1011111011" => n11 <= "10100110111000111010010000011100";
        when "1011111100" => n11 <= "10100110100110111010010001100010";
        when "1011111101" => n11 <= "10100110010100111010010010101001";
        when "1011111110" => n11 <= "10100110000011001010010011101111";
        when "1011111111" => n11 <= "10100101110001001010010100110110";
        when "1100000000" => n11 <= "10100101011111011010010101111101";
        when "1100000001" => n11 <= "10100101001101101010010111000100";
        when "1100000010" => n11 <= "10100100111011111010011000001100";
        when "1100000011" => n11 <= "10100100101010011010011001010011";
        when "1100000100" => n11 <= "10100100011000101010011010011011";
        when "1100000101" => n11 <= "10100100000111001010011011100011";
        when "1100000110" => n11 <= "10100011110101101010011100101011";
        when "1100000111" => n11 <= "10100011100100011010011101110100";
        when "1100001000" => n11 <= "10100011010010111010011110111101";
        when "1100001001" => n11 <= "10100011000001101010100000000110";
        when "1100001010" => n11 <= "10100010110000011010100001001111";
        when "1100001011" => n11 <= "10100010011111001010100010011000";
        when "1100001100" => n11 <= "10100010001110001010100011100010";
        when "1100001101" => n11 <= "10100001111101001010100100101011";
        when "1100001110" => n11 <= "10100001101011111010100101110101";
        when "1100001111" => n11 <= "10100001011011001010100110111111";
        when "1100010000" => n11 <= "10100001001010001010101000001010";
        when "1100010001" => n11 <= "10100000111001011010101001010100";
        when "1100010010" => n11 <= "10100000101000011010101010011111";
        when "1100010011" => n11 <= "10100000010111111010101011101010";
        when "1100010100" => n11 <= "10100000000111001010101100110101";
        when "1100010101" => n11 <= "10011111110110011010101110000001";
        when "1100010110" => n11 <= "10011111100101111010101111001100";
        when "1100010111" => n11 <= "10011111010101011010110000011000";
        when "1100011000" => n11 <= "10011111000100111010110001100100";
        when "1100011001" => n11 <= "10011110110100101010110010110001";
        when "1100011010" => n11 <= "10011110100100001010110011111101";
        when "1100011011" => n11 <= "10011110010011111010110101001010";
        when "1100011100" => n11 <= "10011110000011101010110110010110";
        when "1100011101" => n11 <= "10011101110011101010110111100011";
        when "1100011110" => n11 <= "10011101100011101010111000110001";
        when "1100011111" => n11 <= "10011101010011011010111001111110";
        when "1100100000" => n11 <= "10011101000011011010111011001100";
        when "1100100001" => n11 <= "10011100110011101010111100011010";
        when "1100100010" => n11 <= "10011100100011101010111101101000";
        when "1100100011" => n11 <= "10011100010011111010111110110110";
        when "1100100100" => n11 <= "10011100000100001011000000000100";
        when "1100100101" => n11 <= "10011011110100101011000001010011";
        when "1100100110" => n11 <= "10011011100100111011000010100001";
        when "1100100111" => n11 <= "10011011010101011011000011110000";
        when "1100101000" => n11 <= "10011011000101111011000101000000";
        when "1100101001" => n11 <= "10011010110110011011000110001111";
        when "1100101010" => n11 <= "10011010100111001011000111011110";
        when "1100101011" => n11 <= "10011010010111111011001000101110";
        when "1100101100" => n11 <= "10011010001000101011001001111110";
        when "1100101101" => n11 <= "10011001111001011011001011001110";
        when "1100101110" => n11 <= "10011001101010001011001100011110";
        when "1100101111" => n11 <= "10011001011011001011001101101111";
        when "1100110000" => n11 <= "10011001001100001011001111000000";
        when "1100110001" => n11 <= "10011000111101001011010000010000";
        when "1100110010" => n11 <= "10011000101110011011010001100001";
        when "1100110011" => n11 <= "10011000011111011011010010110011";
        when "1100110100" => n11 <= "10011000010000101011010100000100";
        when "1100110101" => n11 <= "10011000000010001011010101010110";
        when "1100110110" => n11 <= "10010111110011011011010110100111";
        when "1100110111" => n11 <= "10010111100100111011010111111001";
        when "1100111000" => n11 <= "10010111010110011011011001001011";
        when "1100111001" => n11 <= "10010111000111111011011010011110";
        when "1100111010" => n11 <= "10010110111001101011011011110000";
        when "1100111011" => n11 <= "10010110101011001011011101000011";
        when "1100111100" => n11 <= "10010110011100111011011110010110";
        when "1100111101" => n11 <= "10010110001110111011011111101001";
        when "1100111110" => n11 <= "10010110000000101011100000111100";
        when "1100111111" => n11 <= "10010101110010101011100010001111";
        when "1101000000" => n11 <= "10010101100100101011100011100011";
        when "1101000001" => n11 <= "10010101010110101011100100110110";
        when "1101000010" => n11 <= "10010101001000111011100110001010";
        when "1101000011" => n11 <= "10010100111011001011100111011110";
        when "1101000100" => n11 <= "10010100101101011011101000110010";
        when "1101000101" => n11 <= "10010100011111101011101010000111";
        when "1101000110" => n11 <= "10010100010001111011101011011011";
        when "1101000111" => n11 <= "10010100000100011011101100110000";
        when "1101001000" => n11 <= "10010011110110111011101110000101";
        when "1101001001" => n11 <= "10010011101001101011101111011010";
        when "1101001010" => n11 <= "10010011011100001011110000101111";
        when "1101001011" => n11 <= "10010011001110111011110010000100";
        when "1101001100" => n11 <= "10010011000001101011110011011010";
        when "1101001101" => n11 <= "10010010110100101011110100101111";
        when "1101001110" => n11 <= "10010010100111011011110110000101";
        when "1101001111" => n11 <= "10010010011010011011110111011011";
        when "1101010000" => n11 <= "10010010001101011011111000110001";
        when "1101010001" => n11 <= "10010010000000101011111010001000";
        when "1101010010" => n11 <= "10010001110011111011111011011110";
        when "1101010011" => n11 <= "10010001100111001011111100110101";
        when "1101010100" => n11 <= "10010001011010011011111110001100";
        when "1101010101" => n11 <= "10010001001101101011111111100010";
        when "1101010110" => n11 <= "10010001000001001100000000111010";
        when "1101010111" => n11 <= "10010000110100101100000010010001";
        when "1101011000" => n11 <= "10010000101000001100000011101000";
        when "1101011001" => n11 <= "10010000011011111100000101000000";
        when "1101011010" => n11 <= "10010000001111101100000110010111";
        when "1101011011" => n11 <= "10010000000011011100000111101111";
        when "1101011100" => n11 <= "10001111110111001100001001000111";
        when "1101011101" => n11 <= "10001111101011001100001010011111";
        when "1101011110" => n11 <= "10001111011111001100001011111000";
        when "1101011111" => n11 <= "10001111010011001100001101010000";
        when "1101100000" => n11 <= "10001111000111011100001110101001";
        when "1101100001" => n11 <= "10001110111011011100010000000010";
        when "1101100010" => n11 <= "10001110101111101100010001011010";
        when "1101100011" => n11 <= "10001110100100001100010010110011";
        when "1101100100" => n11 <= "10001110011000011100010100001101";
        when "1101100101" => n11 <= "10001110001100111100010101100110";
        when "1101100110" => n11 <= "10001110000001011100010110111111";
        when "1101100111" => n11 <= "10001101110110001100011000011001";
        when "1101101000" => n11 <= "10001101101010101100011001110011";
        when "1101101001" => n11 <= "10001101011111011100011011001101";
        when "1101101010" => n11 <= "10001101010100001100011100100111";
        when "1101101011" => n11 <= "10001101001001001100011110000001";
        when "1101101100" => n11 <= "10001100111110001100011111011011";
        when "1101101101" => n11 <= "10001100110011001100100000110101";
        when "1101101110" => n11 <= "10001100101000001100100010010000";
        when "1101101111" => n11 <= "10001100011101011100100011101011";
        when "1101110000" => n11 <= "10001100010010101100100101000101";
        when "1101110001" => n11 <= "10001100000111111100100110100000";
        when "1101110010" => n11 <= "10001011111101001100100111111011";
        when "1101110011" => n11 <= "10001011110010101100101001010111";
        when "1101110100" => n11 <= "10001011101000001100101010110010";
        when "1101110101" => n11 <= "10001011011101101100101100001101";
        when "1101110110" => n11 <= "10001011010011011100101101101001";
        when "1101110111" => n11 <= "10001011001001001100101111000101";
        when "1101111000" => n11 <= "10001010111110111100110000100001";
        when "1101111001" => n11 <= "10001010110100101100110001111101";
        when "1101111010" => n11 <= "10001010101010101100110011011001";
        when "1101111011" => n11 <= "10001010100000101100110100110101";
        when "1101111100" => n11 <= "10001010010110101100110110010001";
        when "1101111101" => n11 <= "10001010001100111100110111101110";
        when "1101111110" => n11 <= "10001010000010111100111001001010";
        when "1101111111" => n11 <= "10001001111001001100111010100111";
        when "1110000000" => n11 <= "10001001101111101100111100000100";
        when "1110000001" => n11 <= "10001001100101111100111101100001";
        when "1110000010" => n11 <= "10001001011100011100111110111110";
        when "1110000011" => n11 <= "10001001010011001101000000011011";
        when "1110000100" => n11 <= "10001001001001101101000001111000";
        when "1110000101" => n11 <= "10001001000000011101000011010110";
        when "1110000110" => n11 <= "10001000110111001101000100110011";
        when "1110000111" => n11 <= "10001000101110001101000110010001";
        when "1110001000" => n11 <= "10001000100100111101000111101110";
        when "1110001001" => n11 <= "10001000011011111101001001001100";
        when "1110001010" => n11 <= "10001000010010111101001010101010";
        when "1110001011" => n11 <= "10001000001010001101001100001000";
        when "1110001100" => n11 <= "10001000000001011101001101100111";
        when "1110001101" => n11 <= "10000111111000101101001111000101";
        when "1110001110" => n11 <= "10000111101111111101010000100011";
        when "1110001111" => n11 <= "10000111100111011101010010000010";
        when "1110010000" => n11 <= "10000111011110111101010011100000";
        when "1110010001" => n11 <= "10000111010110011101010100111111";
        when "1110010010" => n11 <= "10000111001110001101010110011110";
        when "1110010011" => n11 <= "10000111000101111101010111111101";
        when "1110010100" => n11 <= "10000110111101101101011001011100";
        when "1110010101" => n11 <= "10000110110101011101011010111011";
        when "1110010110" => n11 <= "10000110101101011101011100011010";
        when "1110010111" => n11 <= "10000110100101011101011101111001";
        when "1110011000" => n11 <= "10000110011101011101011111011001";
        when "1110011001" => n11 <= "10000110010101101101100000111000";
        when "1110011010" => n11 <= "10000110001101111101100010011000";
        when "1110011011" => n11 <= "10000110000110001101100011111000";
        when "1110011100" => n11 <= "10000101111110101101100101010111";
        when "1110011101" => n11 <= "10000101110110111101100110110111";
        when "1110011110" => n11 <= "10000101101111011101101000010111";
        when "1110011111" => n11 <= "10000101101000001101101001110111";
        when "1110100000" => n11 <= "10000101100000101101101011010111";
        when "1110100001" => n11 <= "10000101011001011101101100111000";
        when "1110100010" => n11 <= "10000101010010011101101110011000";
        when "1110100011" => n11 <= "10000101001011001101101111111000";
        when "1110100100" => n11 <= "10000101000100001101110001011001";
        when "1110100101" => n11 <= "10000100111101001101110010111010";
        when "1110100110" => n11 <= "10000100110110011101110100011010";
        when "1110100111" => n11 <= "10000100101111011101110101111011";
        when "1110101000" => n11 <= "10000100101000101101110111011100";
        when "1110101001" => n11 <= "10000100100010001101111000111101";
        when "1110101010" => n11 <= "10000100011011011101111010011110";
        when "1110101011" => n11 <= "10000100010100111101111011111111";
        when "1110101100" => n11 <= "10000100001110101101111101100000";
        when "1110101101" => n11 <= "10000100001000001101111111000001";
        when "1110101110" => n11 <= "10000100000001111110000000100011";
        when "1110101111" => n11 <= "10000011111011101110000010000100";
        when "1110110000" => n11 <= "10000011110101101110000011100110";
        when "1110110001" => n11 <= "10000011101111011110000101000111";
        when "1110110010" => n11 <= "10000011101001011110000110101001";
        when "1110110011" => n11 <= "10000011100011101110001000001010";
        when "1110110100" => n11 <= "10000011011101101110001001101100";
        when "1110110101" => n11 <= "10000011010111111110001011001110";
        when "1110110110" => n11 <= "10000011010010001110001100110000";
        when "1110110111" => n11 <= "10000011001100101110001110010010";
        when "1110111000" => n11 <= "10000011000111001110001111110100";
        when "1110111001" => n11 <= "10000011000001101110010001010110";
        when "1110111010" => n11 <= "10000010111100001110010010111000";
        when "1110111011" => n11 <= "10000010110110111110010100011011";
        when "1110111100" => n11 <= "10000010110001101110010101111101";
        when "1110111101" => n11 <= "10000010101100011110010111011111";
        when "1110111110" => n11 <= "10000010100111011110011001000010";
        when "1110111111" => n11 <= "10000010100010011110011010100100";
        when "1111000000" => n11 <= "10000010011101011110011100000111";
        when "1111000001" => n11 <= "10000010011000101110011101101001";
        when "1111000010" => n11 <= "10000010010011111110011111001100";
        when "1111000011" => n11 <= "10000010001111001110100000101111";
        when "1111000100" => n11 <= "10000010001010011110100010010010";
        when "1111000101" => n11 <= "10000010000101111110100011110101";
        when "1111000110" => n11 <= "10000010000001011110100101010111";
        when "1111000111" => n11 <= "10000001111100111110100110111010";
        when "1111001000" => n11 <= "10000001111000101110101000011101";
        when "1111001001" => n11 <= "10000001110100011110101010000000";
        when "1111001010" => n11 <= "10000001110000001110101011100100";
        when "1111001011" => n11 <= "10000001101100001110101101000111";
        when "1111001100" => n11 <= "10000001101000001110101110101010";
        when "1111001101" => n11 <= "10000001100100001110110000001101";
        when "1111001110" => n11 <= "10000001100000001110110001110001";
        when "1111001111" => n11 <= "10000001011100011110110011010100";
        when "1111010000" => n11 <= "10000001011000101110110100110111";
        when "1111010001" => n11 <= "10000001010101001110110110011011";
        when "1111010010" => n11 <= "10000001010001011110110111111110";
        when "1111010011" => n11 <= "10000001001101111110111001100010";
        when "1111010100" => n11 <= "10000001001010101110111011000110";
        when "1111010101" => n11 <= "10000001000111001110111100101001";
        when "1111010110" => n11 <= "10000001000011111110111110001101";
        when "1111010111" => n11 <= "10000001000000101110111111110001";
        when "1111011000" => n11 <= "10000000111101101111000001010100";
        when "1111011001" => n11 <= "10000000111010101111000010111000";
        when "1111011010" => n11 <= "10000000110111101111000100011100";
        when "1111011011" => n11 <= "10000000110100101111000110000000";
        when "1111011100" => n11 <= "10000000110001111111000111100100";
        when "1111011101" => n11 <= "10000000101111001111001001001000";
        when "1111011110" => n11 <= "10000000101100101111001010101100";
        when "1111011111" => n11 <= "10000000101001111111001100010000";
        when "1111100000" => n11 <= "10000000100111011111001101110100";
        when "1111100001" => n11 <= "10000000100101001111001111011000";
        when "1111100010" => n11 <= "10000000100010101111010000111100";
        when "1111100011" => n11 <= "10000000100000011111010010100000";
        when "1111100100" => n11 <= "10000000011110001111010100000100";
        when "1111100101" => n11 <= "10000000011100001111010101101000";
        when "1111100110" => n11 <= "10000000011010001111010111001100";
        when "1111100111" => n11 <= "10000000011000001111011000110001";
        when "1111101000" => n11 <= "10000000010110001111011010010101";
        when "1111101001" => n11 <= "10000000010100011111011011111001";
        when "1111101010" => n11 <= "10000000010010101111011101011101";
        when "1111101011" => n11 <= "10000000010000111111011111000010";
        when "1111101100" => n11 <= "10000000001111011111100000100110";
        when "1111101101" => n11 <= "10000000001101111111100010001010";
        when "1111101110" => n11 <= "10000000001100011111100011101111";
        when "1111101111" => n11 <= "10000000001011001111100101010011";
        when "1111110000" => n11 <= "10000000001001111111100110111000";
        when "1111110001" => n11 <= "10000000001000101111101000011100";
        when "1111110010" => n11 <= "10000000000111101111101010000000";
        when "1111110011" => n11 <= "10000000000110101111101011100101";
        when "1111110100" => n11 <= "10000000000101101111101101001001";
        when "1111110101" => n11 <= "10000000000100101111101110101110";
        when "1111110110" => n11 <= "10000000000011111111110000010010";
        when "1111110111" => n11 <= "10000000000011001111110001110111";
        when "1111111000" => n11 <= "10000000000010011111110011011011";
        when "1111111001" => n11 <= "10000000000001111111110101000000";
        when "1111111010" => n11 <= "10000000000001011111110110100100";
        when "1111111011" => n11 <= "10000000000000111111111000001001";
        when "1111111100" => n11 <= "10000000000000101111111001101101";
        when "1111111101" => n11 <= "10000000000000011111111011010010";
        when "1111111110" => n11 <= "10000000000000001111111100110110";
        when "1111111111" => n11 <= "10000000000000001111111110011011";
        when others => n11 <= "XXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX";
      end case;
    end if;
  end if;
end process;
n12 <= n11(31 downto 31) &
  n11(30 downto 30) &
  n11(29 downto 29) &
  n11(28 downto 28) &
  n11(27 downto 27) &
  n11(26 downto 26) &
  n11(25 downto 25) &
  n11(24 downto 24) &
  n11(23 downto 23) &
  n11(22 downto 22) &
  n11(21 downto 21) &
  n11(20 downto 20) &
  n11(19 downto 19) &
  n11(18 downto 18) &
  n11(17 downto 17) &
  n11(16 downto 16);
n13 <= n11(15 downto 15) &
  n11(14 downto 14) &
  n11(13 downto 13) &
  n11(12 downto 12) &
  n11(11 downto 11) &
  n11(10 downto 10) &
  n11(9 downto 9) &
  n11(8 downto 8) &
  n11(7 downto 7) &
  n11(6 downto 6) &
  n11(5 downto 5) &
  n11(4 downto 4) &
  n11(3 downto 3) &
  n11(2 downto 2) &
  n11(1 downto 1) &
  n11(0 downto 0);
n14 <= unsigned(signed(n5) * signed(n12));
n15 <= n14(30 downto 30) &
  n14(29 downto 29) &
  n14(28 downto 28) &
  n14(27 downto 27) &
  n14(26 downto 26) &
  n14(25 downto 25) &
  n14(24 downto 24) &
  n14(23 downto 23) &
  n14(22 downto 22) &
  n14(21 downto 21) &
  n14(20 downto 20) &
  n14(19 downto 19) &
  n14(18 downto 18) &
  n14(17 downto 17) &
  n14(16 downto 16) &
  n14(15 downto 15);
process (clock_c) begin
  if rising_edge(clock_c) then
    if i5 = "1" then
      n16 <= "0000000000000000";
    elsif i4 = "1" then
      n16 <= n15;
    end if;
  end if;
end process;
n17 <= unsigned(signed(n6) * signed(n13));
n18 <= n17(30 downto 30) &
  n17(29 downto 29) &
  n17(28 downto 28) &
  n17(27 downto 27) &
  n17(26 downto 26) &
  n17(25 downto 25) &
  n17(24 downto 24) &
  n17(23 downto 23) &
  n17(22 downto 22) &
  n17(21 downto 21) &
  n17(20 downto 20) &
  n17(19 downto 19) &
  n17(18 downto 18) &
  n17(17 downto 17) &
  n17(16 downto 16) &
  n17(15 downto 15);
process (clock_c) begin
  if rising_edge(clock_c) then
    if i5 = "1" then
      n19 <= "0000000000000000";
    elsif i4 = "1" then
      n19 <= n18;
    end if;
  end if;
end process;
n20 <= n16 - n19;
process (clock_c) begin
  if rising_edge(clock_c) then
    if i5 = "1" then
      n21 <= "0000000000000000";
    elsif i4 = "1" then
      n21 <= n20;
    end if;
  end if;
end process;
n22 <= unsigned(signed(n5) * signed(n13));
n23 <= n22(30 downto 30) &
  n22(29 downto 29) &
  n22(28 downto 28) &
  n22(27 downto 27) &
  n22(26 downto 26) &
  n22(25 downto 25) &
  n22(24 downto 24) &
  n22(23 downto 23) &
  n22(22 downto 22) &
  n22(21 downto 21) &
  n22(20 downto 20) &
  n22(19 downto 19) &
  n22(18 downto 18) &
  n22(17 downto 17) &
  n22(16 downto 16) &
  n22(15 downto 15);
process (clock_c) begin
  if rising_edge(clock_c) then
    if i5 = "1" then
      n24 <= "0000000000000000";
    elsif i4 = "1" then
      n24 <= n23;
    end if;
  end if;
end process;
n25 <= unsigned(signed(n6) * signed(n12));
n26 <= n25(30 downto 30) &
  n25(29 downto 29) &
  n25(28 downto 28) &
  n25(27 downto 27) &
  n25(26 downto 26) &
  n25(25 downto 25) &
  n25(24 downto 24) &
  n25(23 downto 23) &
  n25(22 downto 22) &
  n25(21 downto 21) &
  n25(20 downto 20) &
  n25(19 downto 19) &
  n25(18 downto 18) &
  n25(17 downto 17) &
  n25(16 downto 16) &
  n25(15 downto 15);
process (clock_c) begin
  if rising_edge(clock_c) then
    if i5 = "1" then
      n27 <= "0000000000000000";
    elsif i4 = "1" then
      n27 <= n26;
    end if;
  end if;
end process;
n28 <= n24 + n27;
process (clock_c) begin
  if rising_edge(clock_c) then
    if i5 = "1" then
      n29 <= "0000000000000000";
    elsif i4 = "1" then
      n29 <= n28;
    end if;
  end if;
end process;
n30 <= n8 + n21;
n31 <= n10 + n29;
n32 <= n30 & n31;
process (clock_c) begin
  if rising_edge(clock_c) then
    if i5 = "1" then
      n33 <= "00000000000000000000000000000000";
    elsif i4 = "1" then
      n33 <= n32;
    end if;
  end if;
end process;
n34 <= n8 - n21;
n35 <= n10 - n29;
n36 <= n34 & n35;
process (clock_c) begin
  if rising_edge(clock_c) then
    if i5 = "1" then
      n37 <= "00000000000000000000000000000000";
    elsif i4 = "1" then
      n37 <= n36;
    end if;
  end if;
end process;
o2 <= n37;
o1 <= n33;
end architecture rtl;

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
entity cf_fft_2048_16_23 is
port (
clock_c : in std_logic;
i1 : in  unsigned(0 downto 0);
i2 : in  unsigned(31 downto 0);
i3 : in  unsigned(31 downto 0);
i4 : in  unsigned(0 downto 0);
i5 : in  unsigned(0 downto 0);
o1 : out unsigned(0 downto 0);
o2 : out unsigned(31 downto 0);
o3 : out unsigned(31 downto 0));
end entity cf_fft_2048_16_23;
architecture rtl of cf_fft_2048_16_23 is
signal n1 : unsigned(9 downto 0);
signal n2 : unsigned(63 downto 0);
signal n3 : unsigned(0 downto 0) := "0";
signal n4 : unsigned(0 downto 0) := "0";
signal n5 : unsigned(0 downto 0) := "0";
signal n6 : unsigned(0 downto 0) := "0";
signal n7 : unsigned(8 downto 0);
signal n8 : unsigned(8 downto 0) := "000000000";
signal n9 : unsigned(8 downto 0) := "000000000";
signal n10 : unsigned(8 downto 0) := "000000000";
signal n11 : unsigned(8 downto 0) := "000000000";
signal n12 : unsigned(0 downto 0);
signal n13 : unsigned(0 downto 0) := "0";
signal n14 : unsigned(0 downto 0) := "0";
signal n15 : unsigned(0 downto 0) := "0";
signal n16 : unsigned(0 downto 0) := "0";
signal n17 : unsigned(0 downto 0);
signal n18 : unsigned(1 downto 0);
signal n19 : unsigned(31 downto 0);
signal n20 : unsigned(31 downto 0);
signal n21 : unsigned(31 downto 0);
signal n22 : unsigned(31 downto 0);
signal n23 : unsigned(31 downto 0);
signal n24 : unsigned(31 downto 0);
signal s25_1 : unsigned(31 downto 0);
signal s25_2 : unsigned(31 downto 0);
signal s26_1 : unsigned(0 downto 0);
signal s27_1 : unsigned(63 downto 0);
signal s28_1 : unsigned(0 downto 0);
signal s28_2 : unsigned(0 downto 0);
signal s28_3 : unsigned(63 downto 0);
signal s29_1 : unsigned(9 downto 0);
signal s29_2 : unsigned(0 downto 0);
component cf_fft_2048_16_24 is
port (
clock_c : in std_logic;
i1 : in  unsigned(31 downto 0);
i2 : in  unsigned(31 downto 0);
i3 : in  unsigned(9 downto 0);
i4 : in  unsigned(0 downto 0);
i5 : in  unsigned(0 downto 0);
o1 : out unsigned(31 downto 0);
o2 : out unsigned(31 downto 0));
end component cf_fft_2048_16_24;
component cf_fft_2048_16_35 is
port (
clock_c : in std_logic;
i1 : in  unsigned(1 downto 0);
i2 : in  unsigned(0 downto 0);
i3 : in  unsigned(0 downto 0);
o1 : out unsigned(0 downto 0));
end component cf_fft_2048_16_35;
component cf_fft_2048_16_31 is
port (
clock_c : in std_logic;
i1 : in  unsigned(63 downto 0);
i2 : in  unsigned(0 downto 0);
i3 : in  unsigned(8 downto 0);
i4 : in  unsigned(0 downto 0);
i5 : in  unsigned(0 downto 0);
i6 : in  unsigned(0 downto 0);
o1 : out unsigned(63 downto 0));
end component cf_fft_2048_16_31;
component cf_fft_2048_16_30 is
port (
clock_c : in std_logic;
i1 : in  unsigned(63 downto 0);
i2 : in  unsigned(0 downto 0);
i3 : in  unsigned(8 downto 0);
i4 : in  unsigned(0 downto 0);
i5 : in  unsigned(0 downto 0);
i6 : in  unsigned(0 downto 0);
o1 : out unsigned(0 downto 0);
o2 : out unsigned(0 downto 0);
o3 : out unsigned(63 downto 0));
end component cf_fft_2048_16_30;
component cf_fft_2048_16_26 is
port (
clock_c : in std_logic;
i1 : in  unsigned(0 downto 0);
i2 : in  unsigned(0 downto 0);
i3 : in  unsigned(0 downto 0);
o1 : out unsigned(9 downto 0);
o2 : out unsigned(0 downto 0));
end component cf_fft_2048_16_26;
begin
n1 <= s29_1(9 downto 9) &
  s29_1(8 downto 8) &
  s29_1(7 downto 7) &
  s29_1(6 downto 6) &
  s29_1(5 downto 5) &
  s29_1(4 downto 4) &
  s29_1(3 downto 3) &
  s29_1(2 downto 2) &
  s29_1(1 downto 1) &
  s29_1(0 downto 0);
n2 <= s25_1 & s25_2;
process (clock_c) begin
  if rising_edge(clock_c) then
    if i5 = "1" then
      n3 <= "0";
    elsif i4 = "1" then
      n3 <= s29_2;
    end if;
  end if;
end process;
process (clock_c) begin
  if rising_edge(clock_c) then
    if i5 = "1" then
      n4 <= "0";
    elsif i4 = "1" then
      n4 <= n3;
    end if;
  end if;
end process;
process (clock_c) begin
  if rising_edge(clock_c) then
    if i5 = "1" then
      n5 <= "0";
    elsif i4 = "1" then
      n5 <= n4;
    end if;
  end if;
end process;
process (clock_c) begin
  if rising_edge(clock_c) then
    if i5 = "1" then
      n6 <= "0";
    elsif i4 = "1" then
      n6 <= n5;
    end if;
  end if;
end process;
n7 <= s29_1(9 downto 9) &
  s29_1(8 downto 8) &
  s29_1(7 downto 7) &
  s29_1(6 downto 6) &
  s29_1(5 downto 5) &
  s29_1(4 downto 4) &
  s29_1(3 downto 3) &
  s29_1(2 downto 2) &
  s29_1(1 downto 1);
process (clock_c) begin
  if rising_edge(clock_c) then
    if i5 = "1" then
      n8 <= "000000000";
    elsif i4 = "1" then
      n8 <= n7;
    end if;
  end if;
end process;
process (clock_c) begin
  if rising_edge(clock_c) then
    if i5 = "1" then
      n9 <= "000000000";
    elsif i4 = "1" then
      n9 <= n8;
    end if;
  end if;
end process;
process (clock_c) begin
  if rising_edge(clock_c) then
    if i5 = "1" then
      n10 <= "000000000";
    elsif i4 = "1" then
      n10 <= n9;
    end if;
  end if;
end process;
process (clock_c) begin
  if rising_edge(clock_c) then
    if i5 = "1" then
      n11 <= "000000000";
    elsif i4 = "1" then
      n11 <= n10;
    end if;
  end if;
end process;
n12 <= s29_1(0 downto 0);
process (clock_c) begin
  if rising_edge(clock_c) then
    if i5 = "1" then
      n13 <= "0";
    elsif i4 = "1" then
      n13 <= n12;
    end if;
  end if;
end process;
process (clock_c) begin
  if rising_edge(clock_c) then
    if i5 = "1" then
      n14 <= "0";
    elsif i4 = "1" then
      n14 <= n13;
    end if;
  end if;
end process;
process (clock_c) begin
  if rising_edge(clock_c) then
    if i5 = "1" then
      n15 <= "0";
    elsif i4 = "1" then
      n15 <= n14;
    end if;
  end if;
end process;
process (clock_c) begin
  if rising_edge(clock_c) then
    if i5 = "1" then
      n16 <= "0";
    elsif i4 = "1" then
      n16 <= n15;
    end if;
  end if;
end process;
n17 <= not n16;
n18 <= s28_2 & s28_1;
n19 <= s28_3(63 downto 63) &
  s28_3(62 downto 62) &
  s28_3(61 downto 61) &
  s28_3(60 downto 60) &
  s28_3(59 downto 59) &
  s28_3(58 downto 58) &
  s28_3(57 downto 57) &
  s28_3(56 downto 56) &
  s28_3(55 downto 55) &
  s28_3(54 downto 54) &
  s28_3(53 downto 53) &
  s28_3(52 downto 52) &
  s28_3(51 downto 51) &
  s28_3(50 downto 50) &
  s28_3(49 downto 49) &
  s28_3(48 downto 48) &
  s28_3(47 downto 47) &
  s28_3(46 downto 46) &
  s28_3(45 downto 45) &
  s28_3(44 downto 44) &
  s28_3(43 downto 43) &
  s28_3(42 downto 42) &
  s28_3(41 downto 41) &
  s28_3(40 downto 40) &
  s28_3(39 downto 39) &
  s28_3(38 downto 38) &
  s28_3(37 downto 37) &
  s28_3(36 downto 36) &
  s28_3(35 downto 35) &
  s28_3(34 downto 34) &
  s28_3(33 downto 33) &
  s28_3(32 downto 32);
n20 <= s28_3(31 downto 31) &
  s28_3(30 downto 30) &
  s28_3(29 downto 29) &
  s28_3(28 downto 28) &
  s28_3(27 downto 27) &
  s28_3(26 downto 26) &
  s28_3(25 downto 25) &
  s28_3(24 downto 24) &
  s28_3(23 downto 23) &
  s28_3(22 downto 22) &
  s28_3(21 downto 21) &
  s28_3(20 downto 20) &
  s28_3(19 downto 19) &
  s28_3(18 downto 18) &
  s28_3(17 downto 17) &
  s28_3(16 downto 16) &
  s28_3(15 downto 15) &
  s28_3(14 downto 14) &
  s28_3(13 downto 13) &
  s28_3(12 downto 12) &
  s28_3(11 downto 11) &
  s28_3(10 downto 10) &
  s28_3(9 downto 9) &
  s28_3(8 downto 8) &
  s28_3(7 downto 7) &
  s28_3(6 downto 6) &
  s28_3(5 downto 5) &
  s28_3(4 downto 4) &
  s28_3(3 downto 3) &
  s28_3(2 downto 2) &
  s28_3(1 downto 1) &
  s28_3(0 downto 0);
n21 <= s27_1(63 downto 63) &
  s27_1(62 downto 62) &
  s27_1(61 downto 61) &
  s27_1(60 downto 60) &
  s27_1(59 downto 59) &
  s27_1(58 downto 58) &
  s27_1(57 downto 57) &
  s27_1(56 downto 56) &
  s27_1(55 downto 55) &
  s27_1(54 downto 54) &
  s27_1(53 downto 53) &
  s27_1(52 downto 52) &
  s27_1(51 downto 51) &
  s27_1(50 downto 50) &
  s27_1(49 downto 49) &
  s27_1(48 downto 48) &
  s27_1(47 downto 47) &
  s27_1(46 downto 46) &
  s27_1(45 downto 45) &
  s27_1(44 downto 44) &
  s27_1(43 downto 43) &
  s27_1(42 downto 42) &
  s27_1(41 downto 41) &
  s27_1(40 downto 40) &
  s27_1(39 downto 39) &
  s27_1(38 downto 38) &
  s27_1(37 downto 37) &
  s27_1(36 downto 36) &
  s27_1(35 downto 35) &
  s27_1(34 downto 34) &
  s27_1(33 downto 33) &
  s27_1(32 downto 32);
n22 <= s27_1(31 downto 31) &
  s27_1(30 downto 30) &
  s27_1(29 downto 29) &
  s27_1(28 downto 28) &
  s27_1(27 downto 27) &
  s27_1(26 downto 26) &
  s27_1(25 downto 25) &
  s27_1(24 downto 24) &
  s27_1(23 downto 23) &
  s27_1(22 downto 22) &
  s27_1(21 downto 21) &
  s27_1(20 downto 20) &
  s27_1(19 downto 19) &
  s27_1(18 downto 18) &
  s27_1(17 downto 17) &
  s27_1(16 downto 16) &
  s27_1(15 downto 15) &
  s27_1(14 downto 14) &
  s27_1(13 downto 13) &
  s27_1(12 downto 12) &
  s27_1(11 downto 11) &
  s27_1(10 downto 10) &
  s27_1(9 downto 9) &
  s27_1(8 downto 8) &
  s27_1(7 downto 7) &
  s27_1(6 downto 6) &
  s27_1(5 downto 5) &
  s27_1(4 downto 4) &
  s27_1(3 downto 3) &
  s27_1(2 downto 2) &
  s27_1(1 downto 1) &
  s27_1(0 downto 0);
n23 <= n20 when s26_1 = "1" else n19;
n24 <= n22 when s26_1 = "1" else n21;
s25 : cf_fft_2048_16_24 port map (clock_c, i2, i3, n1, i4, i5, s25_1, s25_2);
s26 : cf_fft_2048_16_35 port map (clock_c, n18, i4, i5, s26_1);
s27 : cf_fft_2048_16_31 port map (clock_c, n2, n6, n11, n16, i4, i5, s27_1);
s28 : cf_fft_2048_16_30 port map (clock_c, n2, n6, n11, n17, i4, i5, s28_1, s28_2, s28_3);
s29 : cf_fft_2048_16_26 port map (clock_c, i1, i4, i5, s29_1, s29_2);
o3 <= n24;
o2 <= n23;
o1 <= s28_1;
end architecture rtl;

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
entity cf_fft_2048_16_22 is
port (
clock_c : in std_logic;
i1 : in  unsigned(31 downto 0);
i2 : in  unsigned(31 downto 0);
i3 : in  unsigned(8 downto 0);
i4 : in  unsigned(0 downto 0);
i5 : in  unsigned(0 downto 0);
o1 : out unsigned(31 downto 0);
o2 : out unsigned(31 downto 0));
end entity cf_fft_2048_16_22;
architecture rtl of cf_fft_2048_16_22 is
signal n1 : unsigned(31 downto 0) := "00000000000000000000000000000000";
signal n2 : unsigned(15 downto 0);
signal n3 : unsigned(15 downto 0);
signal n4 : unsigned(31 downto 0) := "00000000000000000000000000000000";
signal n5 : unsigned(15 downto 0);
signal n6 : unsigned(15 downto 0);
signal n7 : unsigned(15 downto 0) := "0000000000000000";
signal n8 : unsigned(15 downto 0) := "0000000000000000";
signal n9 : unsigned(15 downto 0) := "0000000000000000";
signal n10 : unsigned(15 downto 0) := "0000000000000000";
signal n11 : unsigned(31 downto 0) := "00000000000000000000000000000000";
signal n12 : unsigned(15 downto 0);
signal n13 : unsigned(15 downto 0);
signal n14 : unsigned(31 downto 0);
signal n15 : unsigned(15 downto 0);
signal n16 : unsigned(15 downto 0) := "0000000000000000";
signal n17 : unsigned(31 downto 0);
signal n18 : unsigned(15 downto 0);
signal n19 : unsigned(15 downto 0) := "0000000000000000";
signal n20 : unsigned(15 downto 0);
signal n21 : unsigned(15 downto 0) := "0000000000000000";
signal n22 : unsigned(31 downto 0);
signal n23 : unsigned(15 downto 0);
signal n24 : unsigned(15 downto 0) := "0000000000000000";
signal n25 : unsigned(31 downto 0);
signal n26 : unsigned(15 downto 0);
signal n27 : unsigned(15 downto 0) := "0000000000000000";
signal n28 : unsigned(15 downto 0);
signal n29 : unsigned(15 downto 0) := "0000000000000000";
signal n30 : unsigned(15 downto 0);
signal n31 : unsigned(15 downto 0);
signal n32 : unsigned(31 downto 0);
signal n33 : unsigned(31 downto 0) := "00000000000000000000000000000000";
signal n34 : unsigned(15 downto 0);
signal n35 : unsigned(15 downto 0);
signal n36 : unsigned(31 downto 0);
signal n37 : unsigned(31 downto 0) := "00000000000000000000000000000000";
begin
process (clock_c) begin
  if rising_edge(clock_c) then
    if i5 = "1" then
      n1 <= "00000000000000000000000000000000";
    elsif i4 = "1" then
      n1 <= i1;
    end if;
  end if;
end process;
n2 <= n1(31 downto 31) &
  n1(30 downto 30) &
  n1(29 downto 29) &
  n1(28 downto 28) &
  n1(27 downto 27) &
  n1(26 downto 26) &
  n1(25 downto 25) &
  n1(24 downto 24) &
  n1(23 downto 23) &
  n1(22 downto 22) &
  n1(21 downto 21) &
  n1(20 downto 20) &
  n1(19 downto 19) &
  n1(18 downto 18) &
  n1(17 downto 17) &
  n1(16 downto 16);
n3 <= n1(15 downto 15) &
  n1(14 downto 14) &
  n1(13 downto 13) &
  n1(12 downto 12) &
  n1(11 downto 11) &
  n1(10 downto 10) &
  n1(9 downto 9) &
  n1(8 downto 8) &
  n1(7 downto 7) &
  n1(6 downto 6) &
  n1(5 downto 5) &
  n1(4 downto 4) &
  n1(3 downto 3) &
  n1(2 downto 2) &
  n1(1 downto 1) &
  n1(0 downto 0);
process (clock_c) begin
  if rising_edge(clock_c) then
    if i5 = "1" then
      n4 <= "00000000000000000000000000000000";
    elsif i4 = "1" then
      n4 <= i2;
    end if;
  end if;
end process;
n5 <= n4(31 downto 31) &
  n4(30 downto 30) &
  n4(29 downto 29) &
  n4(28 downto 28) &
  n4(27 downto 27) &
  n4(26 downto 26) &
  n4(25 downto 25) &
  n4(24 downto 24) &
  n4(23 downto 23) &
  n4(22 downto 22) &
  n4(21 downto 21) &
  n4(20 downto 20) &
  n4(19 downto 19) &
  n4(18 downto 18) &
  n4(17 downto 17) &
  n4(16 downto 16);
n6 <= n4(15 downto 15) &
  n4(14 downto 14) &
  n4(13 downto 13) &
  n4(12 downto 12) &
  n4(11 downto 11) &
  n4(10 downto 10) &
  n4(9 downto 9) &
  n4(8 downto 8) &
  n4(7 downto 7) &
  n4(6 downto 6) &
  n4(5 downto 5) &
  n4(4 downto 4) &
  n4(3 downto 3) &
  n4(2 downto 2) &
  n4(1 downto 1) &
  n4(0 downto 0);
process (clock_c) begin
  if rising_edge(clock_c) then
    if i5 = "1" then
      n7 <= "0000000000000000";
    elsif i4 = "1" then
      n7 <= n2;
    end if;
  end if;
end process;
process (clock_c) begin
  if rising_edge(clock_c) then
    if i5 = "1" then
      n8 <= "0000000000000000";
    elsif i4 = "1" then
      n8 <= n7;
    end if;
  end if;
end process;
process (clock_c) begin
  if rising_edge(clock_c) then
    if i5 = "1" then
      n9 <= "0000000000000000";
    elsif i4 = "1" then
      n9 <= n3;
    end if;
  end if;
end process;
process (clock_c) begin
  if rising_edge(clock_c) then
    if i5 = "1" then
      n10 <= "0000000000000000";
    elsif i4 = "1" then
      n10 <= n9;
    end if;
  end if;
end process;
process (clock_c) begin
  if rising_edge(clock_c) then 
    if i4 = "1" then
      case i3 is
        when "000000000" => n11 <= "01111111111111110000000000000000";
        when "000000001" => n11 <= "01111111111111111111111100110110";
        when "000000010" => n11 <= "01111111111111011111111001101101";
        when "000000011" => n11 <= "01111111111110101111110110100100";
        when "000000100" => n11 <= "01111111111101101111110011011011";
        when "000000101" => n11 <= "01111111111100001111110000010010";
        when "000000110" => n11 <= "01111111111010011111101101001001";
        when "000000111" => n11 <= "01111111111000011111101010000000";
        when "000001000" => n11 <= "01111111110110001111100110111000";
        when "000001001" => n11 <= "01111111110011101111100011101111";
        when "000001010" => n11 <= "01111111110000101111100000100110";
        when "000001011" => n11 <= "01111111101101011111011101011101";
        when "000001100" => n11 <= "01111111101001111111011010010101";
        when "000001101" => n11 <= "01111111100101111111010111001100";
        when "000001110" => n11 <= "01111111100001111111010100000100";
        when "000001111" => n11 <= "01111111011101011111010000111100";
        when "000010000" => n11 <= "01111111011000101111001101110100";
        when "000010001" => n11 <= "01111111010011011111001010101100";
        when "000010010" => n11 <= "01111111001110001111000111100100";
        when "000010011" => n11 <= "01111111001000011111000100011100";
        when "000010100" => n11 <= "01111111000010011111000001010100";
        when "000010101" => n11 <= "01111110111100001110111110001101";
        when "000010110" => n11 <= "01111110110101011110111011000110";
        when "000010111" => n11 <= "01111110101110101110110111111110";
        when "000011000" => n11 <= "01111110100111011110110100110111";
        when "000011001" => n11 <= "01111110011111111110110001110001";
        when "000011010" => n11 <= "01111110010111111110101110101010";
        when "000011011" => n11 <= "01111110001111111110101011100100";
        when "000011100" => n11 <= "01111110000111011110101000011101";
        when "000011101" => n11 <= "01111101111110101110100101010111";
        when "000011110" => n11 <= "01111101110101101110100010010010";
        when "000011111" => n11 <= "01111101101100001110011111001100";
        when "000100000" => n11 <= "01111101100010101110011100000111";
        when "000100001" => n11 <= "01111101011000101110011001000010";
        when "000100010" => n11 <= "01111101001110011110010101111101";
        when "000100011" => n11 <= "01111101000011111110010010111000";
        when "000100100" => n11 <= "01111100111000111110001111110100";
        when "000100101" => n11 <= "01111100101101111110001100110000";
        when "000100110" => n11 <= "01111100100010011110001001101100";
        when "000100111" => n11 <= "01111100010110101110000110101001";
        when "000101000" => n11 <= "01111100001010011110000011100110";
        when "000101001" => n11 <= "01111011111110001110000000100011";
        when "000101010" => n11 <= "01111011110001011101111101100000";
        when "000101011" => n11 <= "01111011100100101101111010011110";
        when "000101100" => n11 <= "01111011010111011101110111011100";
        when "000101101" => n11 <= "01111011001001101101110100011010";
        when "000101110" => n11 <= "01111010111011111101110001011001";
        when "000101111" => n11 <= "01111010101101101101101110011000";
        when "000110000" => n11 <= "01111010011111011101101011010111";
        when "000110001" => n11 <= "01111010010000101101101000010111";
        when "000110010" => n11 <= "01111010000001011101100101010111";
        when "000110011" => n11 <= "01111001110010001101100010011000";
        when "000110100" => n11 <= "01111001100010101101011111011001";
        when "000110101" => n11 <= "01111001010010101101011100011010";
        when "000110110" => n11 <= "01111001000010011101011001011100";
        when "000110111" => n11 <= "01111000110001111101010110011110";
        when "000111000" => n11 <= "01111000100001001101010011100000";
        when "000111001" => n11 <= "01111000010000001101010000100011";
        when "000111010" => n11 <= "01110111111110101101001101100111";
        when "000111011" => n11 <= "01110111101101001101001010101010";
        when "000111100" => n11 <= "01110111011011001101000111101110";
        when "000111101" => n11 <= "01110111001000111101000100110011";
        when "000111110" => n11 <= "01110110110110011101000001111000";
        when "000111111" => n11 <= "01110110100011101100111110111110";
        when "001000000" => n11 <= "01110110010000011100111100000100";
        when "001000001" => n11 <= "01110101111101001100111001001010";
        when "001000010" => n11 <= "01110101101001011100110110010001";
        when "001000011" => n11 <= "01110101010101011100110011011001";
        when "001000100" => n11 <= "01110101000001001100110000100001";
        when "001000101" => n11 <= "01110100101100101100101101101001";
        when "001000110" => n11 <= "01110100010111111100101010110010";
        when "001000111" => n11 <= "01110100000010111100100111111011";
        when "001001000" => n11 <= "01110011101101011100100101000101";
        when "001001001" => n11 <= "01110011010111111100100010010000";
        when "001001010" => n11 <= "01110011000001111100011111011011";
        when "001001011" => n11 <= "01110010101011111100011100100111";
        when "001001100" => n11 <= "01110010010101011100011001110011";
        when "001001101" => n11 <= "01110001111110101100010110111111";
        when "001001110" => n11 <= "01110001100111101100010100001101";
        when "001001111" => n11 <= "01110001010000011100010001011010";
        when "001010000" => n11 <= "01110000111000101100001110101001";
        when "001010001" => n11 <= "01110000100000111100001011111000";
        when "001010010" => n11 <= "01110000001000111100001001000111";
        when "001010011" => n11 <= "01101111110000011100000110010111";
        when "001010100" => n11 <= "01101111010111111100000011101000";
        when "001010101" => n11 <= "01101110111110111100000000111010";
        when "001010110" => n11 <= "01101110100101101011111110001100";
        when "001010111" => n11 <= "01101110001100001011111011011110";
        when "001011000" => n11 <= "01101101110010101011111000110001";
        when "001011001" => n11 <= "01101101011000101011110110000101";
        when "001011010" => n11 <= "01101100111110011011110011011010";
        when "001011011" => n11 <= "01101100100011111011110000101111";
        when "001011100" => n11 <= "01101100001001001011101110000101";
        when "001011101" => n11 <= "01101011101110001011101011011011";
        when "001011110" => n11 <= "01101011010010101011101000110010";
        when "001011111" => n11 <= "01101010110111001011100110001010";
        when "001100000" => n11 <= "01101010011011011011100011100011";
        when "001100001" => n11 <= "01101001111111011011100000111100";
        when "001100010" => n11 <= "01101001100011001011011110010110";
        when "001100011" => n11 <= "01101001000110011011011011110000";
        when "001100100" => n11 <= "01101000101001101011011001001011";
        when "001100101" => n11 <= "01101000001100101011010110100111";
        when "001100110" => n11 <= "01100111101111011011010100000100";
        when "001100111" => n11 <= "01100111010001101011010001100001";
        when "001101000" => n11 <= "01100110110011111011001111000000";
        when "001101001" => n11 <= "01100110010101111011001100011110";
        when "001101010" => n11 <= "01100101110111011011001001111110";
        when "001101011" => n11 <= "01100101011000111011000111011110";
        when "001101100" => n11 <= "01100100111010001011000101000000";
        when "001101101" => n11 <= "01100100011011001011000010100001";
        when "001101110" => n11 <= "01100011111011111011000000000100";
        when "001101111" => n11 <= "01100011011100011010111101101000";
        when "001110000" => n11 <= "01100010111100101010111011001100";
        when "001110001" => n11 <= "01100010011100011010111000110001";
        when "001110010" => n11 <= "01100001111100011010110110010110";
        when "001110011" => n11 <= "01100001011011111010110011111101";
        when "001110100" => n11 <= "01100000111011001010110001100100";
        when "001110101" => n11 <= "01100000011010001010101111001100";
        when "001110110" => n11 <= "01011111111000111010101100110101";
        when "001110111" => n11 <= "01011111010111101010101010011111";
        when "001111000" => n11 <= "01011110110101111010101000001010";
        when "001111001" => n11 <= "01011110010100001010100101110101";
        when "001111010" => n11 <= "01011101110001111010100011100010";
        when "001111011" => n11 <= "01011101001111101010100001001111";
        when "001111100" => n11 <= "01011100101101001010011110111101";
        when "001111101" => n11 <= "01011100001010011010011100101011";
        when "001111110" => n11 <= "01011011100111011010011010011011";
        when "001111111" => n11 <= "01011011000100001010011000001100";
        when "010000000" => n11 <= "01011010100000101010010101111101";
        when "010000001" => n11 <= "01011001111100111010010011101111";
        when "010000010" => n11 <= "01011001011001001010010001100010";
        when "010000011" => n11 <= "01011000110101001010001111010110";
        when "010000100" => n11 <= "01011000010000101010001101001011";
        when "010000101" => n11 <= "01010111101100001010001011000001";
        when "010000110" => n11 <= "01010111000111011010001000111000";
        when "010000111" => n11 <= "01010110100010101010000110101111";
        when "010001000" => n11 <= "01010101111101011010000100101000";
        when "010001001" => n11 <= "01010101011000001010000010100001";
        when "010001010" => n11 <= "01010100110010101010000000011100";
        when "010001011" => n11 <= "01010100001100111001111110010111";
        when "010001100" => n11 <= "01010011100110111001111100010011";
        when "010001101" => n11 <= "01010011000000101001111010010000";
        when "010001110" => n11 <= "01010010011010011001111000001110";
        when "010001111" => n11 <= "01010001110011101001110110001110";
        when "010010000" => n11 <= "01010001001100111001110100001101";
        when "010010001" => n11 <= "01010000100101111001110010001110";
        when "010010010" => n11 <= "01001111111110111001110000010000";
        when "010010011" => n11 <= "01001111010111101001101110010011";
        when "010010100" => n11 <= "01001110101111111001101100010111";
        when "010010101" => n11 <= "01001110001000011001101010011100";
        when "010010110" => n11 <= "01001101100000011001101000100010";
        when "010010111" => n11 <= "01001100111000011001100110101000";
        when "010011000" => n11 <= "01001100001111111001100100110000";
        when "010011001" => n11 <= "01001011100111101001100010111001";
        when "010011010" => n11 <= "01001010111110111001100001000010";
        when "010011011" => n11 <= "01001010010110001001011111001101";
        when "010011100" => n11 <= "01001001101101001001011101011001";
        when "010011101" => n11 <= "01001001000011111001011011100110";
        when "010011110" => n11 <= "01001000011010011001011001110011";
        when "010011111" => n11 <= "01000111110000111001011000000010";
        when "010100000" => n11 <= "01000111000111001001010110010010";
        when "010100001" => n11 <= "01000110011101011001010100100011";
        when "010100010" => n11 <= "01000101110011011001010010110101";
        when "010100011" => n11 <= "01000101001001001001010001000111";
        when "010100100" => n11 <= "01000100011110101001001111011011";
        when "010100101" => n11 <= "01000011110100001001001101110000";
        when "010100110" => n11 <= "01000011001001011001001100000110";
        when "010100111" => n11 <= "01000010011110101001001010011101";
        when "010101000" => n11 <= "01000001110011101001001000110101";
        when "010101001" => n11 <= "01000001001000011001000111001111";
        when "010101010" => n11 <= "01000000011100111001000101101001";
        when "010101011" => n11 <= "00111111110001011001000100000100";
        when "010101100" => n11 <= "00111111000101111001000010100000";
        when "010101101" => n11 <= "00111110011010001001000000111110";
        when "010101110" => n11 <= "00111101101110001000111111011100";
        when "010101111" => n11 <= "00111101000001111000111101111100";
        when "010110000" => n11 <= "00111100010101101000111100011101";
        when "010110001" => n11 <= "00111011101001011000111010111110";
        when "010110010" => n11 <= "00111010111100101000111001100001";
        when "010110011" => n11 <= "00111010010000001000111000000101";
        when "010110100" => n11 <= "00111001100011001000110110101010";
        when "010110101" => n11 <= "00111000110110001000110101010000";
        when "010110110" => n11 <= "00111000001001001000110011111000";
        when "010110111" => n11 <= "00110111011011111000110010100000";
        when "010111000" => n11 <= "00110110101110101000110001001010";
        when "010111001" => n11 <= "00110110000001001000101111110100";
        when "010111010" => n11 <= "00110101010011011000101110100000";
        when "010111011" => n11 <= "00110100100101101000101101001101";
        when "010111100" => n11 <= "00110011110111101000101011111011";
        when "010111101" => n11 <= "00110011001001101000101010101010";
        when "010111110" => n11 <= "00110010011011101000101001011010";
        when "010111111" => n11 <= "00110001101101011000101000001011";
        when "011000000" => n11 <= "00110000111110111000100110111110";
        when "011000001" => n11 <= "00110000010000011000100101110001";
        when "011000010" => n11 <= "00101111100001111000100100100110";
        when "011000011" => n11 <= "00101110110011001000100011011100";
        when "011000100" => n11 <= "00101110000100011000100010010011";
        when "011000101" => n11 <= "00101101010101011000100001001011";
        when "011000110" => n11 <= "00101100100110001000100000000101";
        when "011000111" => n11 <= "00101011110111001000011110111111";
        when "011001000" => n11 <= "00101011000111111000011101111011";
        when "011001001" => n11 <= "00101010011000011000011100111000";
        when "011001010" => n11 <= "00101001101000111000011011110110";
        when "011001011" => n11 <= "00101000111001011000011010110101";
        when "011001100" => n11 <= "00101000001001101000011001110101";
        when "011001101" => n11 <= "00100111011001111000011000110111";
        when "011001110" => n11 <= "00100110101010001000010111111010";
        when "011001111" => n11 <= "00100101111010001000010110111101";
        when "011010000" => n11 <= "00100101001010001000010110000010";
        when "011010001" => n11 <= "00100100011001111000010101001001";
        when "011010010" => n11 <= "00100011101001101000010100010000";
        when "011010011" => n11 <= "00100010111001011000010011011001";
        when "011010100" => n11 <= "00100010001000111000010010100010";
        when "011010101" => n11 <= "00100001011000011000010001101101";
        when "011010110" => n11 <= "00100000100111111000010000111010";
        when "011010111" => n11 <= "00011111110111001000010000000111";
        when "011011000" => n11 <= "00011111000110011000001111010110";
        when "011011001" => n11 <= "00011110010101101000001110100101";
        when "011011010" => n11 <= "00011101100100111000001101110110";
        when "011011011" => n11 <= "00011100110011111000001101001000";
        when "011011100" => n11 <= "00011100000010111000001100011100";
        when "011011101" => n11 <= "00011011010001111000001011110000";
        when "011011110" => n11 <= "00011010100000101000001011000110";
        when "011011111" => n11 <= "00011001101111011000001010011101";
        when "011100000" => n11 <= "00011000111110001000001001110101";
        when "011100001" => n11 <= "00011000001100111000001001001111";
        when "011100010" => n11 <= "00010111011011011000001000101001";
        when "011100011" => n11 <= "00010110101010001000001000000101";
        when "011100100" => n11 <= "00010101111000101000000111100010";
        when "011100101" => n11 <= "00010101000110111000000111000000";
        when "011100110" => n11 <= "00010100010101011000000110100000";
        when "011100111" => n11 <= "00010011100011101000000110000000";
        when "011101000" => n11 <= "00010010110010001000000101100010";
        when "011101001" => n11 <= "00010010000000011000000101000101";
        when "011101010" => n11 <= "00010001001110011000000100101010";
        when "011101011" => n11 <= "00010000011100101000000100001111";
        when "011101100" => n11 <= "00001111101010111000000011110110";
        when "011101101" => n11 <= "00001110111000111000000011011110";
        when "011101110" => n11 <= "00001110000110111000000011000111";
        when "011101111" => n11 <= "00001101010100111000000010110010";
        when "011110000" => n11 <= "00001100100010111000000010011101";
        when "011110001" => n11 <= "00001011110000111000000010001010";
        when "011110010" => n11 <= "00001010111110111000000001111000";
        when "011110011" => n11 <= "00001010001100111000000001101000";
        when "011110100" => n11 <= "00001001011010101000000001011000";
        when "011110101" => n11 <= "00001000101000101000000001001010";
        when "011110110" => n11 <= "00000111110110011000000000111101";
        when "011110111" => n11 <= "00000111000100001000000000110001";
        when "011111000" => n11 <= "00000110010001111000000000100111";
        when "011111001" => n11 <= "00000101011111111000000000011110";
        when "011111010" => n11 <= "00000100101101101000000000010110";
        when "011111011" => n11 <= "00000011111011011000000000001111";
        when "011111100" => n11 <= "00000011001001001000000000001001";
        when "011111101" => n11 <= "00000010010110111000000000000101";
        when "011111110" => n11 <= "00000001100100101000000000000010";
        when "011111111" => n11 <= "00000000110010011000000000000000";
        when "100000000" => n11 <= "00000000000000001000000000000000";
        when "100000001" => n11 <= "11111111001101101000000000000000";
        when "100000010" => n11 <= "11111110011011011000000000000010";
        when "100000011" => n11 <= "11111101101001001000000000000101";
        when "100000100" => n11 <= "11111100110110111000000000001001";
        when "100000101" => n11 <= "11111100000100101000000000001111";
        when "100000110" => n11 <= "11111011010010011000000000010110";
        when "100000111" => n11 <= "11111010100000001000000000011110";
        when "100001000" => n11 <= "11111001101110001000000000100111";
        when "100001001" => n11 <= "11111000111011111000000000110001";
        when "100001010" => n11 <= "11111000001001101000000000111101";
        when "100001011" => n11 <= "11110111010111011000000001001010";
        when "100001100" => n11 <= "11110110100101011000000001011000";
        when "100001101" => n11 <= "11110101110011001000000001101000";
        when "100001110" => n11 <= "11110101000001001000000001111000";
        when "100001111" => n11 <= "11110100001111001000000010001010";
        when "100010000" => n11 <= "11110011011101001000000010011101";
        when "100010001" => n11 <= "11110010101011001000000010110010";
        when "100010010" => n11 <= "11110001111001001000000011000111";
        when "100010011" => n11 <= "11110001000111001000000011011110";
        when "100010100" => n11 <= "11110000010101001000000011110110";
        when "100010101" => n11 <= "11101111100011011000000100001111";
        when "100010110" => n11 <= "11101110110001101000000100101010";
        when "100010111" => n11 <= "11101101111111101000000101000101";
        when "100011000" => n11 <= "11101101001101111000000101100010";
        when "100011001" => n11 <= "11101100011100011000000110000000";
        when "100011010" => n11 <= "11101011101010101000000110100000";
        when "100011011" => n11 <= "11101010111001001000000111000000";
        when "100011100" => n11 <= "11101010000111011000000111100010";
        when "100011101" => n11 <= "11101001010101111000001000000101";
        when "100011110" => n11 <= "11101000100100101000001000101001";
        when "100011111" => n11 <= "11100111110011001000001001001111";
        when "100100000" => n11 <= "11100111000001111000001001110101";
        when "100100001" => n11 <= "11100110010000101000001010011101";
        when "100100010" => n11 <= "11100101011111011000001011000110";
        when "100100011" => n11 <= "11100100101110001000001011110000";
        when "100100100" => n11 <= "11100011111101001000001100011100";
        when "100100101" => n11 <= "11100011001100001000001101001000";
        when "100100110" => n11 <= "11100010011011001000001101110110";
        when "100100111" => n11 <= "11100001101010011000001110100101";
        when "100101000" => n11 <= "11100000111001101000001111010110";
        when "100101001" => n11 <= "11100000001000111000010000000111";
        when "100101010" => n11 <= "11011111011000001000010000111010";
        when "100101011" => n11 <= "11011110100111101000010001101101";
        when "100101100" => n11 <= "11011101110111001000010010100010";
        when "100101101" => n11 <= "11011101000110101000010011011001";
        when "100101110" => n11 <= "11011100010110011000010100010000";
        when "100101111" => n11 <= "11011011100110001000010101001001";
        when "100110000" => n11 <= "11011010110101111000010110000010";
        when "100110001" => n11 <= "11011010000101111000010110111101";
        when "100110010" => n11 <= "11011001010101111000010111111010";
        when "100110011" => n11 <= "11011000100110001000011000110111";
        when "100110100" => n11 <= "11010111110110011000011001110101";
        when "100110101" => n11 <= "11010111000110101000011010110101";
        when "100110110" => n11 <= "11010110010111001000011011110110";
        when "100110111" => n11 <= "11010101100111101000011100111000";
        when "100111000" => n11 <= "11010100111000001000011101111011";
        when "100111001" => n11 <= "11010100001000111000011110111111";
        when "100111010" => n11 <= "11010011011001111000100000000101";
        when "100111011" => n11 <= "11010010101010101000100001001011";
        when "100111100" => n11 <= "11010001111011101000100010010011";
        when "100111101" => n11 <= "11010001001100111000100011011100";
        when "100111110" => n11 <= "11010000011110001000100100100110";
        when "100111111" => n11 <= "11001111101111101000100101110001";
        when "101000000" => n11 <= "11001111000001001000100110111110";
        when "101000001" => n11 <= "11001110010010101000101000001011";
        when "101000010" => n11 <= "11001101100100011000101001011010";
        when "101000011" => n11 <= "11001100110110011000101010101010";
        when "101000100" => n11 <= "11001100001000011000101011111011";
        when "101000101" => n11 <= "11001011011010011000101101001101";
        when "101000110" => n11 <= "11001010101100101000101110100000";
        when "101000111" => n11 <= "11001001111110111000101111110100";
        when "101001000" => n11 <= "11001001010001011000110001001010";
        when "101001001" => n11 <= "11001000100100001000110010100000";
        when "101001010" => n11 <= "11000111110110111000110011111000";
        when "101001011" => n11 <= "11000111001001111000110101010000";
        when "101001100" => n11 <= "11000110011100111000110110101010";
        when "101001101" => n11 <= "11000101101111111000111000000101";
        when "101001110" => n11 <= "11000101000011011000111001100001";
        when "101001111" => n11 <= "11000100010110101000111010111110";
        when "101010000" => n11 <= "11000011101010011000111100011101";
        when "101010001" => n11 <= "11000010111110001000111101111100";
        when "101010010" => n11 <= "11000010010001111000111111011100";
        when "101010011" => n11 <= "11000001100101111001000000111110";
        when "101010100" => n11 <= "11000000111010001001000010100000";
        when "101010101" => n11 <= "11000000001110101001000100000100";
        when "101010110" => n11 <= "10111111100011001001000101101001";
        when "101010111" => n11 <= "10111110110111101001000111001111";
        when "101011000" => n11 <= "10111110001100011001001000110101";
        when "101011001" => n11 <= "10111101100001011001001010011101";
        when "101011010" => n11 <= "10111100110110101001001100000110";
        when "101011011" => n11 <= "10111100001011111001001101110000";
        when "101011100" => n11 <= "10111011100001011001001111011011";
        when "101011101" => n11 <= "10111010110110111001010001000111";
        when "101011110" => n11 <= "10111010001100101001010010110101";
        when "101011111" => n11 <= "10111001100010101001010100100011";
        when "101100000" => n11 <= "10111000111000111001010110010010";
        when "101100001" => n11 <= "10111000001111001001011000000010";
        when "101100010" => n11 <= "10110111100101101001011001110011";
        when "101100011" => n11 <= "10110110111100001001011011100110";
        when "101100100" => n11 <= "10110110010010111001011101011001";
        when "101100101" => n11 <= "10110101101001111001011111001101";
        when "101100110" => n11 <= "10110101000001001001100001000010";
        when "101100111" => n11 <= "10110100011000011001100010111001";
        when "101101000" => n11 <= "10110011110000001001100100110000";
        when "101101001" => n11 <= "10110011000111101001100110101000";
        when "101101010" => n11 <= "10110010011111101001101000100010";
        when "101101011" => n11 <= "10110001110111101001101010011100";
        when "101101100" => n11 <= "10110001010000001001101100010111";
        when "101101101" => n11 <= "10110000101000011001101110010011";
        when "101101110" => n11 <= "10110000000001001001110000010000";
        when "101101111" => n11 <= "10101111011010001001110010001110";
        when "101110000" => n11 <= "10101110110011001001110100001101";
        when "101110001" => n11 <= "10101110001100011001110110001110";
        when "101110010" => n11 <= "10101101100101101001111000001110";
        when "101110011" => n11 <= "10101100111111011001111010010000";
        when "101110100" => n11 <= "10101100011001001001111100010011";
        when "101110101" => n11 <= "10101011110011001001111110010111";
        when "101110110" => n11 <= "10101011001101011010000000011100";
        when "101110111" => n11 <= "10101010100111111010000010100001";
        when "101111000" => n11 <= "10101010000010101010000100101000";
        when "101111001" => n11 <= "10101001011101011010000110101111";
        when "101111010" => n11 <= "10101000111000101010001000111000";
        when "101111011" => n11 <= "10101000010011111010001011000001";
        when "101111100" => n11 <= "10100111101111011010001101001011";
        when "101111101" => n11 <= "10100111001010111010001111010110";
        when "101111110" => n11 <= "10100110100110111010010001100010";
        when "101111111" => n11 <= "10100110000011001010010011101111";
        when "110000000" => n11 <= "10100101011111011010010101111101";
        when "110000001" => n11 <= "10100100111011111010011000001100";
        when "110000010" => n11 <= "10100100011000101010011010011011";
        when "110000011" => n11 <= "10100011110101101010011100101011";
        when "110000100" => n11 <= "10100011010010111010011110111101";
        when "110000101" => n11 <= "10100010110000011010100001001111";
        when "110000110" => n11 <= "10100010001110001010100011100010";
        when "110000111" => n11 <= "10100001101011111010100101110101";
        when "110001000" => n11 <= "10100001001010001010101000001010";
        when "110001001" => n11 <= "10100000101000011010101010011111";
        when "110001010" => n11 <= "10100000000111001010101100110101";
        when "110001011" => n11 <= "10011111100101111010101111001100";
        when "110001100" => n11 <= "10011111000100111010110001100100";
        when "110001101" => n11 <= "10011110100100001010110011111101";
        when "110001110" => n11 <= "10011110000011101010110110010110";
        when "110001111" => n11 <= "10011101100011101010111000110001";
        when "110010000" => n11 <= "10011101000011011010111011001100";
        when "110010001" => n11 <= "10011100100011101010111101101000";
        when "110010010" => n11 <= "10011100000100001011000000000100";
        when "110010011" => n11 <= "10011011100100111011000010100001";
        when "110010100" => n11 <= "10011011000101111011000101000000";
        when "110010101" => n11 <= "10011010100111001011000111011110";
        when "110010110" => n11 <= "10011010001000101011001001111110";
        when "110010111" => n11 <= "10011001101010001011001100011110";
        when "110011000" => n11 <= "10011001001100001011001111000000";
        when "110011001" => n11 <= "10011000101110011011010001100001";
        when "110011010" => n11 <= "10011000010000101011010100000100";
        when "110011011" => n11 <= "10010111110011011011010110100111";
        when "110011100" => n11 <= "10010111010110011011011001001011";
        when "110011101" => n11 <= "10010110111001101011011011110000";
        when "110011110" => n11 <= "10010110011100111011011110010110";
        when "110011111" => n11 <= "10010110000000101011100000111100";
        when "110100000" => n11 <= "10010101100100101011100011100011";
        when "110100001" => n11 <= "10010101001000111011100110001010";
        when "110100010" => n11 <= "10010100101101011011101000110010";
        when "110100011" => n11 <= "10010100010001111011101011011011";
        when "110100100" => n11 <= "10010011110110111011101110000101";
        when "110100101" => n11 <= "10010011011100001011110000101111";
        when "110100110" => n11 <= "10010011000001101011110011011010";
        when "110100111" => n11 <= "10010010100111011011110110000101";
        when "110101000" => n11 <= "10010010001101011011111000110001";
        when "110101001" => n11 <= "10010001110011111011111011011110";
        when "110101010" => n11 <= "10010001011010011011111110001100";
        when "110101011" => n11 <= "10010001000001001100000000111010";
        when "110101100" => n11 <= "10010000101000001100000011101000";
        when "110101101" => n11 <= "10010000001111101100000110010111";
        when "110101110" => n11 <= "10001111110111001100001001000111";
        when "110101111" => n11 <= "10001111011111001100001011111000";
        when "110110000" => n11 <= "10001111000111011100001110101001";
        when "110110001" => n11 <= "10001110101111101100010001011010";
        when "110110010" => n11 <= "10001110011000011100010100001101";
        when "110110011" => n11 <= "10001110000001011100010110111111";
        when "110110100" => n11 <= "10001101101010101100011001110011";
        when "110110101" => n11 <= "10001101010100001100011100100111";
        when "110110110" => n11 <= "10001100111110001100011111011011";
        when "110110111" => n11 <= "10001100101000001100100010010000";
        when "110111000" => n11 <= "10001100010010101100100101000101";
        when "110111001" => n11 <= "10001011111101001100100111111011";
        when "110111010" => n11 <= "10001011101000001100101010110010";
        when "110111011" => n11 <= "10001011010011011100101101101001";
        when "110111100" => n11 <= "10001010111110111100110000100001";
        when "110111101" => n11 <= "10001010101010101100110011011001";
        when "110111110" => n11 <= "10001010010110101100110110010001";
        when "110111111" => n11 <= "10001010000010111100111001001010";
        when "111000000" => n11 <= "10001001101111101100111100000100";
        when "111000001" => n11 <= "10001001011100011100111110111110";
        when "111000010" => n11 <= "10001001001001101101000001111000";
        when "111000011" => n11 <= "10001000110111001101000100110011";
        when "111000100" => n11 <= "10001000100100111101000111101110";
        when "111000101" => n11 <= "10001000010010111101001010101010";
        when "111000110" => n11 <= "10001000000001011101001101100111";
        when "111000111" => n11 <= "10000111101111111101010000100011";
        when "111001000" => n11 <= "10000111011110111101010011100000";
        when "111001001" => n11 <= "10000111001110001101010110011110";
        when "111001010" => n11 <= "10000110111101101101011001011100";
        when "111001011" => n11 <= "10000110101101011101011100011010";
        when "111001100" => n11 <= "10000110011101011101011111011001";
        when "111001101" => n11 <= "10000110001101111101100010011000";
        when "111001110" => n11 <= "10000101111110101101100101010111";
        when "111001111" => n11 <= "10000101101111011101101000010111";
        when "111010000" => n11 <= "10000101100000101101101011010111";
        when "111010001" => n11 <= "10000101010010011101101110011000";
        when "111010010" => n11 <= "10000101000100001101110001011001";
        when "111010011" => n11 <= "10000100110110011101110100011010";
        when "111010100" => n11 <= "10000100101000101101110111011100";
        when "111010101" => n11 <= "10000100011011011101111010011110";
        when "111010110" => n11 <= "10000100001110101101111101100000";
        when "111010111" => n11 <= "10000100000001111110000000100011";
        when "111011000" => n11 <= "10000011110101101110000011100110";
        when "111011001" => n11 <= "10000011101001011110000110101001";
        when "111011010" => n11 <= "10000011011101101110001001101100";
        when "111011011" => n11 <= "10000011010010001110001100110000";
        when "111011100" => n11 <= "10000011000111001110001111110100";
        when "111011101" => n11 <= "10000010111100001110010010111000";
        when "111011110" => n11 <= "10000010110001101110010101111101";
        when "111011111" => n11 <= "10000010100111011110011001000010";
        when "111100000" => n11 <= "10000010011101011110011100000111";
        when "111100001" => n11 <= "10000010010011111110011111001100";
        when "111100010" => n11 <= "10000010001010011110100010010010";
        when "111100011" => n11 <= "10000010000001011110100101010111";
        when "111100100" => n11 <= "10000001111000101110101000011101";
        when "111100101" => n11 <= "10000001110000001110101011100100";
        when "111100110" => n11 <= "10000001101000001110101110101010";
        when "111100111" => n11 <= "10000001100000001110110001110001";
        when "111101000" => n11 <= "10000001011000101110110100110111";
        when "111101001" => n11 <= "10000001010001011110110111111110";
        when "111101010" => n11 <= "10000001001010101110111011000110";
        when "111101011" => n11 <= "10000001000011111110111110001101";
        when "111101100" => n11 <= "10000000111101101111000001010100";
        when "111101101" => n11 <= "10000000110111101111000100011100";
        when "111101110" => n11 <= "10000000110001111111000111100100";
        when "111101111" => n11 <= "10000000101100101111001010101100";
        when "111110000" => n11 <= "10000000100111011111001101110100";
        when "111110001" => n11 <= "10000000100010101111010000111100";
        when "111110010" => n11 <= "10000000011110001111010100000100";
        when "111110011" => n11 <= "10000000011010001111010111001100";
        when "111110100" => n11 <= "10000000010110001111011010010101";
        when "111110101" => n11 <= "10000000010010101111011101011101";
        when "111110110" => n11 <= "10000000001111011111100000100110";
        when "111110111" => n11 <= "10000000001100011111100011101111";
        when "111111000" => n11 <= "10000000001001111111100110111000";
        when "111111001" => n11 <= "10000000000111101111101010000000";
        when "111111010" => n11 <= "10000000000101101111101101001001";
        when "111111011" => n11 <= "10000000000011111111110000010010";
        when "111111100" => n11 <= "10000000000010011111110011011011";
        when "111111101" => n11 <= "10000000000001011111110110100100";
        when "111111110" => n11 <= "10000000000000101111111001101101";
        when "111111111" => n11 <= "10000000000000001111111100110110";
        when others => n11 <= "XXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX";
      end case;
    end if;
  end if;
end process;
n12 <= n11(31 downto 31) &
  n11(30 downto 30) &
  n11(29 downto 29) &
  n11(28 downto 28) &
  n11(27 downto 27) &
  n11(26 downto 26) &
  n11(25 downto 25) &
  n11(24 downto 24) &
  n11(23 downto 23) &
  n11(22 downto 22) &
  n11(21 downto 21) &
  n11(20 downto 20) &
  n11(19 downto 19) &
  n11(18 downto 18) &
  n11(17 downto 17) &
  n11(16 downto 16);
n13 <= n11(15 downto 15) &
  n11(14 downto 14) &
  n11(13 downto 13) &
  n11(12 downto 12) &
  n11(11 downto 11) &
  n11(10 downto 10) &
  n11(9 downto 9) &
  n11(8 downto 8) &
  n11(7 downto 7) &
  n11(6 downto 6) &
  n11(5 downto 5) &
  n11(4 downto 4) &
  n11(3 downto 3) &
  n11(2 downto 2) &
  n11(1 downto 1) &
  n11(0 downto 0);
n14 <= unsigned(signed(n5) * signed(n12));
n15 <= n14(30 downto 30) &
  n14(29 downto 29) &
  n14(28 downto 28) &
  n14(27 downto 27) &
  n14(26 downto 26) &
  n14(25 downto 25) &
  n14(24 downto 24) &
  n14(23 downto 23) &
  n14(22 downto 22) &
  n14(21 downto 21) &
  n14(20 downto 20) &
  n14(19 downto 19) &
  n14(18 downto 18) &
  n14(17 downto 17) &
  n14(16 downto 16) &
  n14(15 downto 15);
process (clock_c) begin
  if rising_edge(clock_c) then
    if i5 = "1" then
      n16 <= "0000000000000000";
    elsif i4 = "1" then
      n16 <= n15;
    end if;
  end if;
end process;
n17 <= unsigned(signed(n6) * signed(n13));
n18 <= n17(30 downto 30) &
  n17(29 downto 29) &
  n17(28 downto 28) &
  n17(27 downto 27) &
  n17(26 downto 26) &
  n17(25 downto 25) &
  n17(24 downto 24) &
  n17(23 downto 23) &
  n17(22 downto 22) &
  n17(21 downto 21) &
  n17(20 downto 20) &
  n17(19 downto 19) &
  n17(18 downto 18) &
  n17(17 downto 17) &
  n17(16 downto 16) &
  n17(15 downto 15);
process (clock_c) begin
  if rising_edge(clock_c) then
    if i5 = "1" then
      n19 <= "0000000000000000";
    elsif i4 = "1" then
      n19 <= n18;
    end if;
  end if;
end process;
n20 <= n16 - n19;
process (clock_c) begin
  if rising_edge(clock_c) then
    if i5 = "1" then
      n21 <= "0000000000000000";
    elsif i4 = "1" then
      n21 <= n20;
    end if;
  end if;
end process;
n22 <= unsigned(signed(n5) * signed(n13));
n23 <= n22(30 downto 30) &
  n22(29 downto 29) &
  n22(28 downto 28) &
  n22(27 downto 27) &
  n22(26 downto 26) &
  n22(25 downto 25) &
  n22(24 downto 24) &
  n22(23 downto 23) &
  n22(22 downto 22) &
  n22(21 downto 21) &
  n22(20 downto 20) &
  n22(19 downto 19) &
  n22(18 downto 18) &
  n22(17 downto 17) &
  n22(16 downto 16) &
  n22(15 downto 15);
process (clock_c) begin
  if rising_edge(clock_c) then
    if i5 = "1" then
      n24 <= "0000000000000000";
    elsif i4 = "1" then
      n24 <= n23;
    end if;
  end if;
end process;
n25 <= unsigned(signed(n6) * signed(n12));
n26 <= n25(30 downto 30) &
  n25(29 downto 29) &
  n25(28 downto 28) &
  n25(27 downto 27) &
  n25(26 downto 26) &
  n25(25 downto 25) &
  n25(24 downto 24) &
  n25(23 downto 23) &
  n25(22 downto 22) &
  n25(21 downto 21) &
  n25(20 downto 20) &
  n25(19 downto 19) &
  n25(18 downto 18) &
  n25(17 downto 17) &
  n25(16 downto 16) &
  n25(15 downto 15);
process (clock_c) begin
  if rising_edge(clock_c) then
    if i5 = "1" then
      n27 <= "0000000000000000";
    elsif i4 = "1" then
      n27 <= n26;
    end if;
  end if;
end process;
n28 <= n24 + n27;
process (clock_c) begin
  if rising_edge(clock_c) then
    if i5 = "1" then
      n29 <= "0000000000000000";
    elsif i4 = "1" then
      n29 <= n28;
    end if;
  end if;
end process;
n30 <= n8 + n21;
n31 <= n10 + n29;
n32 <= n30 & n31;
process (clock_c) begin
  if rising_edge(clock_c) then
    if i5 = "1" then
      n33 <= "00000000000000000000000000000000";
    elsif i4 = "1" then
      n33 <= n32;
    end if;
  end if;
end process;
n34 <= n8 - n21;
n35 <= n10 - n29;
n36 <= n34 & n35;
process (clock_c) begin
  if rising_edge(clock_c) then
    if i5 = "1" then
      n37 <= "00000000000000000000000000000000";
    elsif i4 = "1" then
      n37 <= n36;
    end if;
  end if;
end process;
o2 <= n37;
o1 <= n33;
end architecture rtl;

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
entity cf_fft_2048_16_21 is
port (
clock_c : in std_logic;
i1 : in  unsigned(0 downto 0);
i2 : in  unsigned(31 downto 0);
i3 : in  unsigned(31 downto 0);
i4 : in  unsigned(0 downto 0);
i5 : in  unsigned(0 downto 0);
o1 : out unsigned(0 downto 0);
o2 : out unsigned(31 downto 0);
o3 : out unsigned(31 downto 0));
end entity cf_fft_2048_16_21;
architecture rtl of cf_fft_2048_16_21 is
signal n1 : unsigned(8 downto 0);
signal n2 : unsigned(63 downto 0);
signal n3 : unsigned(0 downto 0) := "0";
signal n4 : unsigned(0 downto 0) := "0";
signal n5 : unsigned(0 downto 0) := "0";
signal n6 : unsigned(0 downto 0) := "0";
signal n7 : unsigned(8 downto 0);
signal n8 : unsigned(8 downto 0) := "000000000";
signal n9 : unsigned(8 downto 0) := "000000000";
signal n10 : unsigned(8 downto 0) := "000000000";
signal n11 : unsigned(8 downto 0) := "000000000";
signal n12 : unsigned(0 downto 0);
signal n13 : unsigned(0 downto 0) := "0";
signal n14 : unsigned(0 downto 0) := "0";
signal n15 : unsigned(0 downto 0) := "0";
signal n16 : unsigned(0 downto 0) := "0";
signal n17 : unsigned(0 downto 0);
signal n18 : unsigned(1 downto 0);
signal n19 : unsigned(31 downto 0);
signal n20 : unsigned(31 downto 0);
signal n21 : unsigned(31 downto 0);
signal n22 : unsigned(31 downto 0);
signal n23 : unsigned(31 downto 0);
signal n24 : unsigned(31 downto 0);
signal s25_1 : unsigned(31 downto 0);
signal s25_2 : unsigned(31 downto 0);
signal s26_1 : unsigned(0 downto 0);
signal s27_1 : unsigned(63 downto 0);
signal s28_1 : unsigned(0 downto 0);
signal s28_2 : unsigned(0 downto 0);
signal s28_3 : unsigned(63 downto 0);
signal s29_1 : unsigned(9 downto 0);
signal s29_2 : unsigned(0 downto 0);
component cf_fft_2048_16_22 is
port (
clock_c : in std_logic;
i1 : in  unsigned(31 downto 0);
i2 : in  unsigned(31 downto 0);
i3 : in  unsigned(8 downto 0);
i4 : in  unsigned(0 downto 0);
i5 : in  unsigned(0 downto 0);
o1 : out unsigned(31 downto 0);
o2 : out unsigned(31 downto 0));
end component cf_fft_2048_16_22;
component cf_fft_2048_16_35 is
port (
clock_c : in std_logic;
i1 : in  unsigned(1 downto 0);
i2 : in  unsigned(0 downto 0);
i3 : in  unsigned(0 downto 0);
o1 : out unsigned(0 downto 0));
end component cf_fft_2048_16_35;
component cf_fft_2048_16_31 is
port (
clock_c : in std_logic;
i1 : in  unsigned(63 downto 0);
i2 : in  unsigned(0 downto 0);
i3 : in  unsigned(8 downto 0);
i4 : in  unsigned(0 downto 0);
i5 : in  unsigned(0 downto 0);
i6 : in  unsigned(0 downto 0);
o1 : out unsigned(63 downto 0));
end component cf_fft_2048_16_31;
component cf_fft_2048_16_30 is
port (
clock_c : in std_logic;
i1 : in  unsigned(63 downto 0);
i2 : in  unsigned(0 downto 0);
i3 : in  unsigned(8 downto 0);
i4 : in  unsigned(0 downto 0);
i5 : in  unsigned(0 downto 0);
i6 : in  unsigned(0 downto 0);
o1 : out unsigned(0 downto 0);
o2 : out unsigned(0 downto 0);
o3 : out unsigned(63 downto 0));
end component cf_fft_2048_16_30;
component cf_fft_2048_16_26 is
port (
clock_c : in std_logic;
i1 : in  unsigned(0 downto 0);
i2 : in  unsigned(0 downto 0);
i3 : in  unsigned(0 downto 0);
o1 : out unsigned(9 downto 0);
o2 : out unsigned(0 downto 0));
end component cf_fft_2048_16_26;
begin
n1 <= s29_1(9 downto 9) &
  s29_1(8 downto 8) &
  s29_1(7 downto 7) &
  s29_1(6 downto 6) &
  s29_1(5 downto 5) &
  s29_1(4 downto 4) &
  s29_1(3 downto 3) &
  s29_1(2 downto 2) &
  s29_1(1 downto 1);
n2 <= s25_1 & s25_2;
process (clock_c) begin
  if rising_edge(clock_c) then
    if i5 = "1" then
      n3 <= "0";
    elsif i4 = "1" then
      n3 <= s29_2;
    end if;
  end if;
end process;
process (clock_c) begin
  if rising_edge(clock_c) then
    if i5 = "1" then
      n4 <= "0";
    elsif i4 = "1" then
      n4 <= n3;
    end if;
  end if;
end process;
process (clock_c) begin
  if rising_edge(clock_c) then
    if i5 = "1" then
      n5 <= "0";
    elsif i4 = "1" then
      n5 <= n4;
    end if;
  end if;
end process;
process (clock_c) begin
  if rising_edge(clock_c) then
    if i5 = "1" then
      n6 <= "0";
    elsif i4 = "1" then
      n6 <= n5;
    end if;
  end if;
end process;
n7 <= s29_1(9 downto 9) &
  s29_1(8 downto 8) &
  s29_1(7 downto 7) &
  s29_1(6 downto 6) &
  s29_1(5 downto 5) &
  s29_1(4 downto 4) &
  s29_1(3 downto 3) &
  s29_1(2 downto 2) &
  s29_1(1 downto 1);
process (clock_c) begin
  if rising_edge(clock_c) then
    if i5 = "1" then
      n8 <= "000000000";
    elsif i4 = "1" then
      n8 <= n7;
    end if;
  end if;
end process;
process (clock_c) begin
  if rising_edge(clock_c) then
    if i5 = "1" then
      n9 <= "000000000";
    elsif i4 = "1" then
      n9 <= n8;
    end if;
  end if;
end process;
process (clock_c) begin
  if rising_edge(clock_c) then
    if i5 = "1" then
      n10 <= "000000000";
    elsif i4 = "1" then
      n10 <= n9;
    end if;
  end if;
end process;
process (clock_c) begin
  if rising_edge(clock_c) then
    if i5 = "1" then
      n11 <= "000000000";
    elsif i4 = "1" then
      n11 <= n10;
    end if;
  end if;
end process;
n12 <= s29_1(0 downto 0);
process (clock_c) begin
  if rising_edge(clock_c) then
    if i5 = "1" then
      n13 <= "0";
    elsif i4 = "1" then
      n13 <= n12;
    end if;
  end if;
end process;
process (clock_c) begin
  if rising_edge(clock_c) then
    if i5 = "1" then
      n14 <= "0";
    elsif i4 = "1" then
      n14 <= n13;
    end if;
  end if;
end process;
process (clock_c) begin
  if rising_edge(clock_c) then
    if i5 = "1" then
      n15 <= "0";
    elsif i4 = "1" then
      n15 <= n14;
    end if;
  end if;
end process;
process (clock_c) begin
  if rising_edge(clock_c) then
    if i5 = "1" then
      n16 <= "0";
    elsif i4 = "1" then
      n16 <= n15;
    end if;
  end if;
end process;
n17 <= not n16;
n18 <= s28_2 & s28_1;
n19 <= s28_3(63 downto 63) &
  s28_3(62 downto 62) &
  s28_3(61 downto 61) &
  s28_3(60 downto 60) &
  s28_3(59 downto 59) &
  s28_3(58 downto 58) &
  s28_3(57 downto 57) &
  s28_3(56 downto 56) &
  s28_3(55 downto 55) &
  s28_3(54 downto 54) &
  s28_3(53 downto 53) &
  s28_3(52 downto 52) &
  s28_3(51 downto 51) &
  s28_3(50 downto 50) &
  s28_3(49 downto 49) &
  s28_3(48 downto 48) &
  s28_3(47 downto 47) &
  s28_3(46 downto 46) &
  s28_3(45 downto 45) &
  s28_3(44 downto 44) &
  s28_3(43 downto 43) &
  s28_3(42 downto 42) &
  s28_3(41 downto 41) &
  s28_3(40 downto 40) &
  s28_3(39 downto 39) &
  s28_3(38 downto 38) &
  s28_3(37 downto 37) &
  s28_3(36 downto 36) &
  s28_3(35 downto 35) &
  s28_3(34 downto 34) &
  s28_3(33 downto 33) &
  s28_3(32 downto 32);
n20 <= s28_3(31 downto 31) &
  s28_3(30 downto 30) &
  s28_3(29 downto 29) &
  s28_3(28 downto 28) &
  s28_3(27 downto 27) &
  s28_3(26 downto 26) &
  s28_3(25 downto 25) &
  s28_3(24 downto 24) &
  s28_3(23 downto 23) &
  s28_3(22 downto 22) &
  s28_3(21 downto 21) &
  s28_3(20 downto 20) &
  s28_3(19 downto 19) &
  s28_3(18 downto 18) &
  s28_3(17 downto 17) &
  s28_3(16 downto 16) &
  s28_3(15 downto 15) &
  s28_3(14 downto 14) &
  s28_3(13 downto 13) &
  s28_3(12 downto 12) &
  s28_3(11 downto 11) &
  s28_3(10 downto 10) &
  s28_3(9 downto 9) &
  s28_3(8 downto 8) &
  s28_3(7 downto 7) &
  s28_3(6 downto 6) &
  s28_3(5 downto 5) &
  s28_3(4 downto 4) &
  s28_3(3 downto 3) &
  s28_3(2 downto 2) &
  s28_3(1 downto 1) &
  s28_3(0 downto 0);
n21 <= s27_1(63 downto 63) &
  s27_1(62 downto 62) &
  s27_1(61 downto 61) &
  s27_1(60 downto 60) &
  s27_1(59 downto 59) &
  s27_1(58 downto 58) &
  s27_1(57 downto 57) &
  s27_1(56 downto 56) &
  s27_1(55 downto 55) &
  s27_1(54 downto 54) &
  s27_1(53 downto 53) &
  s27_1(52 downto 52) &
  s27_1(51 downto 51) &
  s27_1(50 downto 50) &
  s27_1(49 downto 49) &
  s27_1(48 downto 48) &
  s27_1(47 downto 47) &
  s27_1(46 downto 46) &
  s27_1(45 downto 45) &
  s27_1(44 downto 44) &
  s27_1(43 downto 43) &
  s27_1(42 downto 42) &
  s27_1(41 downto 41) &
  s27_1(40 downto 40) &
  s27_1(39 downto 39) &
  s27_1(38 downto 38) &
  s27_1(37 downto 37) &
  s27_1(36 downto 36) &
  s27_1(35 downto 35) &
  s27_1(34 downto 34) &
  s27_1(33 downto 33) &
  s27_1(32 downto 32);
n22 <= s27_1(31 downto 31) &
  s27_1(30 downto 30) &
  s27_1(29 downto 29) &
  s27_1(28 downto 28) &
  s27_1(27 downto 27) &
  s27_1(26 downto 26) &
  s27_1(25 downto 25) &
  s27_1(24 downto 24) &
  s27_1(23 downto 23) &
  s27_1(22 downto 22) &
  s27_1(21 downto 21) &
  s27_1(20 downto 20) &
  s27_1(19 downto 19) &
  s27_1(18 downto 18) &
  s27_1(17 downto 17) &
  s27_1(16 downto 16) &
  s27_1(15 downto 15) &
  s27_1(14 downto 14) &
  s27_1(13 downto 13) &
  s27_1(12 downto 12) &
  s27_1(11 downto 11) &
  s27_1(10 downto 10) &
  s27_1(9 downto 9) &
  s27_1(8 downto 8) &
  s27_1(7 downto 7) &
  s27_1(6 downto 6) &
  s27_1(5 downto 5) &
  s27_1(4 downto 4) &
  s27_1(3 downto 3) &
  s27_1(2 downto 2) &
  s27_1(1 downto 1) &
  s27_1(0 downto 0);
n23 <= n20 when s26_1 = "1" else n19;
n24 <= n22 when s26_1 = "1" else n21;
s25 : cf_fft_2048_16_22 port map (clock_c, i2, i3, n1, i4, i5, s25_1, s25_2);
s26 : cf_fft_2048_16_35 port map (clock_c, n18, i4, i5, s26_1);
s27 : cf_fft_2048_16_31 port map (clock_c, n2, n6, n11, n16, i4, i5, s27_1);
s28 : cf_fft_2048_16_30 port map (clock_c, n2, n6, n11, n17, i4, i5, s28_1, s28_2, s28_3);
s29 : cf_fft_2048_16_26 port map (clock_c, i1, i4, i5, s29_1, s29_2);
o3 <= n24;
o2 <= n23;
o1 <= s28_1;
end architecture rtl;

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
entity cf_fft_2048_16_20 is
port (
clock_c : in std_logic;
i1 : in  unsigned(31 downto 0);
i2 : in  unsigned(31 downto 0);
i3 : in  unsigned(7 downto 0);
i4 : in  unsigned(0 downto 0);
i5 : in  unsigned(0 downto 0);
o1 : out unsigned(31 downto 0);
o2 : out unsigned(31 downto 0));
end entity cf_fft_2048_16_20;
architecture rtl of cf_fft_2048_16_20 is
signal n1 : unsigned(31 downto 0) := "00000000000000000000000000000000";
signal n2 : unsigned(15 downto 0);
signal n3 : unsigned(15 downto 0);
signal n4 : unsigned(31 downto 0) := "00000000000000000000000000000000";
signal n5 : unsigned(15 downto 0);
signal n6 : unsigned(15 downto 0);
signal n7 : unsigned(15 downto 0) := "0000000000000000";
signal n8 : unsigned(15 downto 0) := "0000000000000000";
signal n9 : unsigned(15 downto 0) := "0000000000000000";
signal n10 : unsigned(15 downto 0) := "0000000000000000";
signal n11 : unsigned(31 downto 0) := "00000000000000000000000000000000";
signal n12 : unsigned(15 downto 0);
signal n13 : unsigned(15 downto 0);
signal n14 : unsigned(31 downto 0);
signal n15 : unsigned(15 downto 0);
signal n16 : unsigned(15 downto 0) := "0000000000000000";
signal n17 : unsigned(31 downto 0);
signal n18 : unsigned(15 downto 0);
signal n19 : unsigned(15 downto 0) := "0000000000000000";
signal n20 : unsigned(15 downto 0);
signal n21 : unsigned(15 downto 0) := "0000000000000000";
signal n22 : unsigned(31 downto 0);
signal n23 : unsigned(15 downto 0);
signal n24 : unsigned(15 downto 0) := "0000000000000000";
signal n25 : unsigned(31 downto 0);
signal n26 : unsigned(15 downto 0);
signal n27 : unsigned(15 downto 0) := "0000000000000000";
signal n28 : unsigned(15 downto 0);
signal n29 : unsigned(15 downto 0) := "0000000000000000";
signal n30 : unsigned(15 downto 0);
signal n31 : unsigned(15 downto 0);
signal n32 : unsigned(31 downto 0);
signal n33 : unsigned(31 downto 0) := "00000000000000000000000000000000";
signal n34 : unsigned(15 downto 0);
signal n35 : unsigned(15 downto 0);
signal n36 : unsigned(31 downto 0);
signal n37 : unsigned(31 downto 0) := "00000000000000000000000000000000";
begin
process (clock_c) begin
  if rising_edge(clock_c) then
    if i5 = "1" then
      n1 <= "00000000000000000000000000000000";
    elsif i4 = "1" then
      n1 <= i1;
    end if;
  end if;
end process;
n2 <= n1(31 downto 31) &
  n1(30 downto 30) &
  n1(29 downto 29) &
  n1(28 downto 28) &
  n1(27 downto 27) &
  n1(26 downto 26) &
  n1(25 downto 25) &
  n1(24 downto 24) &
  n1(23 downto 23) &
  n1(22 downto 22) &
  n1(21 downto 21) &
  n1(20 downto 20) &
  n1(19 downto 19) &
  n1(18 downto 18) &
  n1(17 downto 17) &
  n1(16 downto 16);
n3 <= n1(15 downto 15) &
  n1(14 downto 14) &
  n1(13 downto 13) &
  n1(12 downto 12) &
  n1(11 downto 11) &
  n1(10 downto 10) &
  n1(9 downto 9) &
  n1(8 downto 8) &
  n1(7 downto 7) &
  n1(6 downto 6) &
  n1(5 downto 5) &
  n1(4 downto 4) &
  n1(3 downto 3) &
  n1(2 downto 2) &
  n1(1 downto 1) &
  n1(0 downto 0);
process (clock_c) begin
  if rising_edge(clock_c) then
    if i5 = "1" then
      n4 <= "00000000000000000000000000000000";
    elsif i4 = "1" then
      n4 <= i2;
    end if;
  end if;
end process;
n5 <= n4(31 downto 31) &
  n4(30 downto 30) &
  n4(29 downto 29) &
  n4(28 downto 28) &
  n4(27 downto 27) &
  n4(26 downto 26) &
  n4(25 downto 25) &
  n4(24 downto 24) &
  n4(23 downto 23) &
  n4(22 downto 22) &
  n4(21 downto 21) &
  n4(20 downto 20) &
  n4(19 downto 19) &
  n4(18 downto 18) &
  n4(17 downto 17) &
  n4(16 downto 16);
n6 <= n4(15 downto 15) &
  n4(14 downto 14) &
  n4(13 downto 13) &
  n4(12 downto 12) &
  n4(11 downto 11) &
  n4(10 downto 10) &
  n4(9 downto 9) &
  n4(8 downto 8) &
  n4(7 downto 7) &
  n4(6 downto 6) &
  n4(5 downto 5) &
  n4(4 downto 4) &
  n4(3 downto 3) &
  n4(2 downto 2) &
  n4(1 downto 1) &
  n4(0 downto 0);
process (clock_c) begin
  if rising_edge(clock_c) then
    if i5 = "1" then
      n7 <= "0000000000000000";
    elsif i4 = "1" then
      n7 <= n2;
    end if;
  end if;
end process;
process (clock_c) begin
  if rising_edge(clock_c) then
    if i5 = "1" then
      n8 <= "0000000000000000";
    elsif i4 = "1" then
      n8 <= n7;
    end if;
  end if;
end process;
process (clock_c) begin
  if rising_edge(clock_c) then
    if i5 = "1" then
      n9 <= "0000000000000000";
    elsif i4 = "1" then
      n9 <= n3;
    end if;
  end if;
end process;
process (clock_c) begin
  if rising_edge(clock_c) then
    if i5 = "1" then
      n10 <= "0000000000000000";
    elsif i4 = "1" then
      n10 <= n9;
    end if;
  end if;
end process;
process (clock_c) begin
  if rising_edge(clock_c) then 
    if i4 = "1" then
      case i3 is
        when "00000000" => n11 <= "01111111111111110000000000000000";
        when "00000001" => n11 <= "01111111111111011111111001101101";
        when "00000010" => n11 <= "01111111111101101111110011011011";
        when "00000011" => n11 <= "01111111111010011111101101001001";
        when "00000100" => n11 <= "01111111110110001111100110111000";
        when "00000101" => n11 <= "01111111110000101111100000100110";
        when "00000110" => n11 <= "01111111101001111111011010010101";
        when "00000111" => n11 <= "01111111100001111111010100000100";
        when "00001000" => n11 <= "01111111011000101111001101110100";
        when "00001001" => n11 <= "01111111001110001111000111100100";
        when "00001010" => n11 <= "01111111000010011111000001010100";
        when "00001011" => n11 <= "01111110110101011110111011000110";
        when "00001100" => n11 <= "01111110100111011110110100110111";
        when "00001101" => n11 <= "01111110010111111110101110101010";
        when "00001110" => n11 <= "01111110000111011110101000011101";
        when "00001111" => n11 <= "01111101110101101110100010010010";
        when "00010000" => n11 <= "01111101100010101110011100000111";
        when "00010001" => n11 <= "01111101001110011110010101111101";
        when "00010010" => n11 <= "01111100111000111110001111110100";
        when "00010011" => n11 <= "01111100100010011110001001101100";
        when "00010100" => n11 <= "01111100001010011110000011100110";
        when "00010101" => n11 <= "01111011110001011101111101100000";
        when "00010110" => n11 <= "01111011010111011101110111011100";
        when "00010111" => n11 <= "01111010111011111101110001011001";
        when "00011000" => n11 <= "01111010011111011101101011010111";
        when "00011001" => n11 <= "01111010000001011101100101010111";
        when "00011010" => n11 <= "01111001100010101101011111011001";
        when "00011011" => n11 <= "01111001000010011101011001011100";
        when "00011100" => n11 <= "01111000100001001101010011100000";
        when "00011101" => n11 <= "01110111111110101101001101100111";
        when "00011110" => n11 <= "01110111011011001101000111101110";
        when "00011111" => n11 <= "01110110110110011101000001111000";
        when "00100000" => n11 <= "01110110010000011100111100000100";
        when "00100001" => n11 <= "01110101101001011100110110010001";
        when "00100010" => n11 <= "01110101000001001100110000100001";
        when "00100011" => n11 <= "01110100010111111100101010110010";
        when "00100100" => n11 <= "01110011101101011100100101000101";
        when "00100101" => n11 <= "01110011000001111100011111011011";
        when "00100110" => n11 <= "01110010010101011100011001110011";
        when "00100111" => n11 <= "01110001100111101100010100001101";
        when "00101000" => n11 <= "01110000111000101100001110101001";
        when "00101001" => n11 <= "01110000001000111100001001000111";
        when "00101010" => n11 <= "01101111010111111100000011101000";
        when "00101011" => n11 <= "01101110100101101011111110001100";
        when "00101100" => n11 <= "01101101110010101011111000110001";
        when "00101101" => n11 <= "01101100111110011011110011011010";
        when "00101110" => n11 <= "01101100001001001011101110000101";
        when "00101111" => n11 <= "01101011010010101011101000110010";
        when "00110000" => n11 <= "01101010011011011011100011100011";
        when "00110001" => n11 <= "01101001100011001011011110010110";
        when "00110010" => n11 <= "01101000101001101011011001001011";
        when "00110011" => n11 <= "01100111101111011011010100000100";
        when "00110100" => n11 <= "01100110110011111011001111000000";
        when "00110101" => n11 <= "01100101110111011011001001111110";
        when "00110110" => n11 <= "01100100111010001011000101000000";
        when "00110111" => n11 <= "01100011111011111011000000000100";
        when "00111000" => n11 <= "01100010111100101010111011001100";
        when "00111001" => n11 <= "01100001111100011010110110010110";
        when "00111010" => n11 <= "01100000111011001010110001100100";
        when "00111011" => n11 <= "01011111111000111010101100110101";
        when "00111100" => n11 <= "01011110110101111010101000001010";
        when "00111101" => n11 <= "01011101110001111010100011100010";
        when "00111110" => n11 <= "01011100101101001010011110111101";
        when "00111111" => n11 <= "01011011100111011010011010011011";
        when "01000000" => n11 <= "01011010100000101010010101111101";
        when "01000001" => n11 <= "01011001011001001010010001100010";
        when "01000010" => n11 <= "01011000010000101010001101001011";
        when "01000011" => n11 <= "01010111000111011010001000111000";
        when "01000100" => n11 <= "01010101111101011010000100101000";
        when "01000101" => n11 <= "01010100110010101010000000011100";
        when "01000110" => n11 <= "01010011100110111001111100010011";
        when "01000111" => n11 <= "01010010011010011001111000001110";
        when "01001000" => n11 <= "01010001001100111001110100001101";
        when "01001001" => n11 <= "01001111111110111001110000010000";
        when "01001010" => n11 <= "01001110101111111001101100010111";
        when "01001011" => n11 <= "01001101100000011001101000100010";
        when "01001100" => n11 <= "01001100001111111001100100110000";
        when "01001101" => n11 <= "01001010111110111001100001000010";
        when "01001110" => n11 <= "01001001101101001001011101011001";
        when "01001111" => n11 <= "01001000011010011001011001110011";
        when "01010000" => n11 <= "01000111000111001001010110010010";
        when "01010001" => n11 <= "01000101110011011001010010110101";
        when "01010010" => n11 <= "01000100011110101001001111011011";
        when "01010011" => n11 <= "01000011001001011001001100000110";
        when "01010100" => n11 <= "01000001110011101001001000110101";
        when "01010101" => n11 <= "01000000011100111001000101101001";
        when "01010110" => n11 <= "00111111000101111001000010100000";
        when "01010111" => n11 <= "00111101101110001000111111011100";
        when "01011000" => n11 <= "00111100010101101000111100011101";
        when "01011001" => n11 <= "00111010111100101000111001100001";
        when "01011010" => n11 <= "00111001100011001000110110101010";
        when "01011011" => n11 <= "00111000001001001000110011111000";
        when "01011100" => n11 <= "00110110101110101000110001001010";
        when "01011101" => n11 <= "00110101010011011000101110100000";
        when "01011110" => n11 <= "00110011110111101000101011111011";
        when "01011111" => n11 <= "00110010011011101000101001011010";
        when "01100000" => n11 <= "00110000111110111000100110111110";
        when "01100001" => n11 <= "00101111100001111000100100100110";
        when "01100010" => n11 <= "00101110000100011000100010010011";
        when "01100011" => n11 <= "00101100100110001000100000000101";
        when "01100100" => n11 <= "00101011000111111000011101111011";
        when "01100101" => n11 <= "00101001101000111000011011110110";
        when "01100110" => n11 <= "00101000001001101000011001110101";
        when "01100111" => n11 <= "00100110101010001000010111111010";
        when "01101000" => n11 <= "00100101001010001000010110000010";
        when "01101001" => n11 <= "00100011101001101000010100010000";
        when "01101010" => n11 <= "00100010001000111000010010100010";
        when "01101011" => n11 <= "00100000100111111000010000111010";
        when "01101100" => n11 <= "00011111000110011000001111010110";
        when "01101101" => n11 <= "00011101100100111000001101110110";
        when "01101110" => n11 <= "00011100000010111000001100011100";
        when "01101111" => n11 <= "00011010100000101000001011000110";
        when "01110000" => n11 <= "00011000111110001000001001110101";
        when "01110001" => n11 <= "00010111011011011000001000101001";
        when "01110010" => n11 <= "00010101111000101000000111100010";
        when "01110011" => n11 <= "00010100010101011000000110100000";
        when "01110100" => n11 <= "00010010110010001000000101100010";
        when "01110101" => n11 <= "00010001001110011000000100101010";
        when "01110110" => n11 <= "00001111101010111000000011110110";
        when "01110111" => n11 <= "00001110000110111000000011000111";
        when "01111000" => n11 <= "00001100100010111000000010011101";
        when "01111001" => n11 <= "00001010111110111000000001111000";
        when "01111010" => n11 <= "00001001011010101000000001011000";
        when "01111011" => n11 <= "00000111110110011000000000111101";
        when "01111100" => n11 <= "00000110010001111000000000100111";
        when "01111101" => n11 <= "00000100101101101000000000010110";
        when "01111110" => n11 <= "00000011001001001000000000001001";
        when "01111111" => n11 <= "00000001100100101000000000000010";
        when "10000000" => n11 <= "00000000000000001000000000000000";
        when "10000001" => n11 <= "11111110011011011000000000000010";
        when "10000010" => n11 <= "11111100110110111000000000001001";
        when "10000011" => n11 <= "11111011010010011000000000010110";
        when "10000100" => n11 <= "11111001101110001000000000100111";
        when "10000101" => n11 <= "11111000001001101000000000111101";
        when "10000110" => n11 <= "11110110100101011000000001011000";
        when "10000111" => n11 <= "11110101000001001000000001111000";
        when "10001000" => n11 <= "11110011011101001000000010011101";
        when "10001001" => n11 <= "11110001111001001000000011000111";
        when "10001010" => n11 <= "11110000010101001000000011110110";
        when "10001011" => n11 <= "11101110110001101000000100101010";
        when "10001100" => n11 <= "11101101001101111000000101100010";
        when "10001101" => n11 <= "11101011101010101000000110100000";
        when "10001110" => n11 <= "11101010000111011000000111100010";
        when "10001111" => n11 <= "11101000100100101000001000101001";
        when "10010000" => n11 <= "11100111000001111000001001110101";
        when "10010001" => n11 <= "11100101011111011000001011000110";
        when "10010010" => n11 <= "11100011111101001000001100011100";
        when "10010011" => n11 <= "11100010011011001000001101110110";
        when "10010100" => n11 <= "11100000111001101000001111010110";
        when "10010101" => n11 <= "11011111011000001000010000111010";
        when "10010110" => n11 <= "11011101110111001000010010100010";
        when "10010111" => n11 <= "11011100010110011000010100010000";
        when "10011000" => n11 <= "11011010110101111000010110000010";
        when "10011001" => n11 <= "11011001010101111000010111111010";
        when "10011010" => n11 <= "11010111110110011000011001110101";
        when "10011011" => n11 <= "11010110010111001000011011110110";
        when "10011100" => n11 <= "11010100111000001000011101111011";
        when "10011101" => n11 <= "11010011011001111000100000000101";
        when "10011110" => n11 <= "11010001111011101000100010010011";
        when "10011111" => n11 <= "11010000011110001000100100100110";
        when "10100000" => n11 <= "11001111000001001000100110111110";
        when "10100001" => n11 <= "11001101100100011000101001011010";
        when "10100010" => n11 <= "11001100001000011000101011111011";
        when "10100011" => n11 <= "11001010101100101000101110100000";
        when "10100100" => n11 <= "11001001010001011000110001001010";
        when "10100101" => n11 <= "11000111110110111000110011111000";
        when "10100110" => n11 <= "11000110011100111000110110101010";
        when "10100111" => n11 <= "11000101000011011000111001100001";
        when "10101000" => n11 <= "11000011101010011000111100011101";
        when "10101001" => n11 <= "11000010010001111000111111011100";
        when "10101010" => n11 <= "11000000111010001001000010100000";
        when "10101011" => n11 <= "10111111100011001001000101101001";
        when "10101100" => n11 <= "10111110001100011001001000110101";
        when "10101101" => n11 <= "10111100110110101001001100000110";
        when "10101110" => n11 <= "10111011100001011001001111011011";
        when "10101111" => n11 <= "10111010001100101001010010110101";
        when "10110000" => n11 <= "10111000111000111001010110010010";
        when "10110001" => n11 <= "10110111100101101001011001110011";
        when "10110010" => n11 <= "10110110010010111001011101011001";
        when "10110011" => n11 <= "10110101000001001001100001000010";
        when "10110100" => n11 <= "10110011110000001001100100110000";
        when "10110101" => n11 <= "10110010011111101001101000100010";
        when "10110110" => n11 <= "10110001010000001001101100010111";
        when "10110111" => n11 <= "10110000000001001001110000010000";
        when "10111000" => n11 <= "10101110110011001001110100001101";
        when "10111001" => n11 <= "10101101100101101001111000001110";
        when "10111010" => n11 <= "10101100011001001001111100010011";
        when "10111011" => n11 <= "10101011001101011010000000011100";
        when "10111100" => n11 <= "10101010000010101010000100101000";
        when "10111101" => n11 <= "10101000111000101010001000111000";
        when "10111110" => n11 <= "10100111101111011010001101001011";
        when "10111111" => n11 <= "10100110100110111010010001100010";
        when "11000000" => n11 <= "10100101011111011010010101111101";
        when "11000001" => n11 <= "10100100011000101010011010011011";
        when "11000010" => n11 <= "10100011010010111010011110111101";
        when "11000011" => n11 <= "10100010001110001010100011100010";
        when "11000100" => n11 <= "10100001001010001010101000001010";
        when "11000101" => n11 <= "10100000000111001010101100110101";
        when "11000110" => n11 <= "10011111000100111010110001100100";
        when "11000111" => n11 <= "10011110000011101010110110010110";
        when "11001000" => n11 <= "10011101000011011010111011001100";
        when "11001001" => n11 <= "10011100000100001011000000000100";
        when "11001010" => n11 <= "10011011000101111011000101000000";
        when "11001011" => n11 <= "10011010001000101011001001111110";
        when "11001100" => n11 <= "10011001001100001011001111000000";
        when "11001101" => n11 <= "10011000010000101011010100000100";
        when "11001110" => n11 <= "10010111010110011011011001001011";
        when "11001111" => n11 <= "10010110011100111011011110010110";
        when "11010000" => n11 <= "10010101100100101011100011100011";
        when "11010001" => n11 <= "10010100101101011011101000110010";
        when "11010010" => n11 <= "10010011110110111011101110000101";
        when "11010011" => n11 <= "10010011000001101011110011011010";
        when "11010100" => n11 <= "10010010001101011011111000110001";
        when "11010101" => n11 <= "10010001011010011011111110001100";
        when "11010110" => n11 <= "10010000101000001100000011101000";
        when "11010111" => n11 <= "10001111110111001100001001000111";
        when "11011000" => n11 <= "10001111000111011100001110101001";
        when "11011001" => n11 <= "10001110011000011100010100001101";
        when "11011010" => n11 <= "10001101101010101100011001110011";
        when "11011011" => n11 <= "10001100111110001100011111011011";
        when "11011100" => n11 <= "10001100010010101100100101000101";
        when "11011101" => n11 <= "10001011101000001100101010110010";
        when "11011110" => n11 <= "10001010111110111100110000100001";
        when "11011111" => n11 <= "10001010010110101100110110010001";
        when "11100000" => n11 <= "10001001101111101100111100000100";
        when "11100001" => n11 <= "10001001001001101101000001111000";
        when "11100010" => n11 <= "10001000100100111101000111101110";
        when "11100011" => n11 <= "10001000000001011101001101100111";
        when "11100100" => n11 <= "10000111011110111101010011100000";
        when "11100101" => n11 <= "10000110111101101101011001011100";
        when "11100110" => n11 <= "10000110011101011101011111011001";
        when "11100111" => n11 <= "10000101111110101101100101010111";
        when "11101000" => n11 <= "10000101100000101101101011010111";
        when "11101001" => n11 <= "10000101000100001101110001011001";
        when "11101010" => n11 <= "10000100101000101101110111011100";
        when "11101011" => n11 <= "10000100001110101101111101100000";
        when "11101100" => n11 <= "10000011110101101110000011100110";
        when "11101101" => n11 <= "10000011011101101110001001101100";
        when "11101110" => n11 <= "10000011000111001110001111110100";
        when "11101111" => n11 <= "10000010110001101110010101111101";
        when "11110000" => n11 <= "10000010011101011110011100000111";
        when "11110001" => n11 <= "10000010001010011110100010010010";
        when "11110010" => n11 <= "10000001111000101110101000011101";
        when "11110011" => n11 <= "10000001101000001110101110101010";
        when "11110100" => n11 <= "10000001011000101110110100110111";
        when "11110101" => n11 <= "10000001001010101110111011000110";
        when "11110110" => n11 <= "10000000111101101111000001010100";
        when "11110111" => n11 <= "10000000110001111111000111100100";
        when "11111000" => n11 <= "10000000100111011111001101110100";
        when "11111001" => n11 <= "10000000011110001111010100000100";
        when "11111010" => n11 <= "10000000010110001111011010010101";
        when "11111011" => n11 <= "10000000001111011111100000100110";
        when "11111100" => n11 <= "10000000001001111111100110111000";
        when "11111101" => n11 <= "10000000000101101111101101001001";
        when "11111110" => n11 <= "10000000000010011111110011011011";
        when "11111111" => n11 <= "10000000000000101111111001101101";
        when others => n11 <= "XXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX";
      end case;
    end if;
  end if;
end process;
n12 <= n11(31 downto 31) &
  n11(30 downto 30) &
  n11(29 downto 29) &
  n11(28 downto 28) &
  n11(27 downto 27) &
  n11(26 downto 26) &
  n11(25 downto 25) &
  n11(24 downto 24) &
  n11(23 downto 23) &
  n11(22 downto 22) &
  n11(21 downto 21) &
  n11(20 downto 20) &
  n11(19 downto 19) &
  n11(18 downto 18) &
  n11(17 downto 17) &
  n11(16 downto 16);
n13 <= n11(15 downto 15) &
  n11(14 downto 14) &
  n11(13 downto 13) &
  n11(12 downto 12) &
  n11(11 downto 11) &
  n11(10 downto 10) &
  n11(9 downto 9) &
  n11(8 downto 8) &
  n11(7 downto 7) &
  n11(6 downto 6) &
  n11(5 downto 5) &
  n11(4 downto 4) &
  n11(3 downto 3) &
  n11(2 downto 2) &
  n11(1 downto 1) &
  n11(0 downto 0);
n14 <= unsigned(signed(n5) * signed(n12));
n15 <= n14(30 downto 30) &
  n14(29 downto 29) &
  n14(28 downto 28) &
  n14(27 downto 27) &
  n14(26 downto 26) &
  n14(25 downto 25) &
  n14(24 downto 24) &
  n14(23 downto 23) &
  n14(22 downto 22) &
  n14(21 downto 21) &
  n14(20 downto 20) &
  n14(19 downto 19) &
  n14(18 downto 18) &
  n14(17 downto 17) &
  n14(16 downto 16) &
  n14(15 downto 15);
process (clock_c) begin
  if rising_edge(clock_c) then
    if i5 = "1" then
      n16 <= "0000000000000000";
    elsif i4 = "1" then
      n16 <= n15;
    end if;
  end if;
end process;
n17 <= unsigned(signed(n6) * signed(n13));
n18 <= n17(30 downto 30) &
  n17(29 downto 29) &
  n17(28 downto 28) &
  n17(27 downto 27) &
  n17(26 downto 26) &
  n17(25 downto 25) &
  n17(24 downto 24) &
  n17(23 downto 23) &
  n17(22 downto 22) &
  n17(21 downto 21) &
  n17(20 downto 20) &
  n17(19 downto 19) &
  n17(18 downto 18) &
  n17(17 downto 17) &
  n17(16 downto 16) &
  n17(15 downto 15);
process (clock_c) begin
  if rising_edge(clock_c) then
    if i5 = "1" then
      n19 <= "0000000000000000";
    elsif i4 = "1" then
      n19 <= n18;
    end if;
  end if;
end process;
n20 <= n16 - n19;
process (clock_c) begin
  if rising_edge(clock_c) then
    if i5 = "1" then
      n21 <= "0000000000000000";
    elsif i4 = "1" then
      n21 <= n20;
    end if;
  end if;
end process;
n22 <= unsigned(signed(n5) * signed(n13));
n23 <= n22(30 downto 30) &
  n22(29 downto 29) &
  n22(28 downto 28) &
  n22(27 downto 27) &
  n22(26 downto 26) &
  n22(25 downto 25) &
  n22(24 downto 24) &
  n22(23 downto 23) &
  n22(22 downto 22) &
  n22(21 downto 21) &
  n22(20 downto 20) &
  n22(19 downto 19) &
  n22(18 downto 18) &
  n22(17 downto 17) &
  n22(16 downto 16) &
  n22(15 downto 15);
process (clock_c) begin
  if rising_edge(clock_c) then
    if i5 = "1" then
      n24 <= "0000000000000000";
    elsif i4 = "1" then
      n24 <= n23;
    end if;
  end if;
end process;
n25 <= unsigned(signed(n6) * signed(n12));
n26 <= n25(30 downto 30) &
  n25(29 downto 29) &
  n25(28 downto 28) &
  n25(27 downto 27) &
  n25(26 downto 26) &
  n25(25 downto 25) &
  n25(24 downto 24) &
  n25(23 downto 23) &
  n25(22 downto 22) &
  n25(21 downto 21) &
  n25(20 downto 20) &
  n25(19 downto 19) &
  n25(18 downto 18) &
  n25(17 downto 17) &
  n25(16 downto 16) &
  n25(15 downto 15);
process (clock_c) begin
  if rising_edge(clock_c) then
    if i5 = "1" then
      n27 <= "0000000000000000";
    elsif i4 = "1" then
      n27 <= n26;
    end if;
  end if;
end process;
n28 <= n24 + n27;
process (clock_c) begin
  if rising_edge(clock_c) then
    if i5 = "1" then
      n29 <= "0000000000000000";
    elsif i4 = "1" then
      n29 <= n28;
    end if;
  end if;
end process;
n30 <= n8 + n21;
n31 <= n10 + n29;
n32 <= n30 & n31;
process (clock_c) begin
  if rising_edge(clock_c) then
    if i5 = "1" then
      n33 <= "00000000000000000000000000000000";
    elsif i4 = "1" then
      n33 <= n32;
    end if;
  end if;
end process;
n34 <= n8 - n21;
n35 <= n10 - n29;
n36 <= n34 & n35;
process (clock_c) begin
  if rising_edge(clock_c) then
    if i5 = "1" then
      n37 <= "00000000000000000000000000000000";
    elsif i4 = "1" then
      n37 <= n36;
    end if;
  end if;
end process;
o2 <= n37;
o1 <= n33;
end architecture rtl;

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
entity cf_fft_2048_16_19 is
port (
clock_c : in std_logic;
i1 : in  unsigned(0 downto 0);
i2 : in  unsigned(31 downto 0);
i3 : in  unsigned(31 downto 0);
i4 : in  unsigned(0 downto 0);
i5 : in  unsigned(0 downto 0);
o1 : out unsigned(0 downto 0);
o2 : out unsigned(31 downto 0);
o3 : out unsigned(31 downto 0));
end entity cf_fft_2048_16_19;
architecture rtl of cf_fft_2048_16_19 is
signal n1 : unsigned(7 downto 0);
signal n2 : unsigned(63 downto 0);
signal n3 : unsigned(0 downto 0) := "0";
signal n4 : unsigned(0 downto 0) := "0";
signal n5 : unsigned(0 downto 0) := "0";
signal n6 : unsigned(0 downto 0) := "0";
signal n7 : unsigned(8 downto 0);
signal n8 : unsigned(8 downto 0) := "000000000";
signal n9 : unsigned(8 downto 0) := "000000000";
signal n10 : unsigned(8 downto 0) := "000000000";
signal n11 : unsigned(8 downto 0) := "000000000";
signal n12 : unsigned(0 downto 0);
signal n13 : unsigned(0 downto 0) := "0";
signal n14 : unsigned(0 downto 0) := "0";
signal n15 : unsigned(0 downto 0) := "0";
signal n16 : unsigned(0 downto 0) := "0";
signal n17 : unsigned(0 downto 0);
signal n18 : unsigned(1 downto 0);
signal n19 : unsigned(31 downto 0);
signal n20 : unsigned(31 downto 0);
signal n21 : unsigned(31 downto 0);
signal n22 : unsigned(31 downto 0);
signal n23 : unsigned(31 downto 0);
signal n24 : unsigned(31 downto 0);
signal s25_1 : unsigned(31 downto 0);
signal s25_2 : unsigned(31 downto 0);
signal s26_1 : unsigned(0 downto 0);
signal s27_1 : unsigned(63 downto 0);
signal s28_1 : unsigned(0 downto 0);
signal s28_2 : unsigned(0 downto 0);
signal s28_3 : unsigned(63 downto 0);
signal s29_1 : unsigned(9 downto 0);
signal s29_2 : unsigned(0 downto 0);
component cf_fft_2048_16_20 is
port (
clock_c : in std_logic;
i1 : in  unsigned(31 downto 0);
i2 : in  unsigned(31 downto 0);
i3 : in  unsigned(7 downto 0);
i4 : in  unsigned(0 downto 0);
i5 : in  unsigned(0 downto 0);
o1 : out unsigned(31 downto 0);
o2 : out unsigned(31 downto 0));
end component cf_fft_2048_16_20;
component cf_fft_2048_16_35 is
port (
clock_c : in std_logic;
i1 : in  unsigned(1 downto 0);
i2 : in  unsigned(0 downto 0);
i3 : in  unsigned(0 downto 0);
o1 : out unsigned(0 downto 0));
end component cf_fft_2048_16_35;
component cf_fft_2048_16_31 is
port (
clock_c : in std_logic;
i1 : in  unsigned(63 downto 0);
i2 : in  unsigned(0 downto 0);
i3 : in  unsigned(8 downto 0);
i4 : in  unsigned(0 downto 0);
i5 : in  unsigned(0 downto 0);
i6 : in  unsigned(0 downto 0);
o1 : out unsigned(63 downto 0));
end component cf_fft_2048_16_31;
component cf_fft_2048_16_30 is
port (
clock_c : in std_logic;
i1 : in  unsigned(63 downto 0);
i2 : in  unsigned(0 downto 0);
i3 : in  unsigned(8 downto 0);
i4 : in  unsigned(0 downto 0);
i5 : in  unsigned(0 downto 0);
i6 : in  unsigned(0 downto 0);
o1 : out unsigned(0 downto 0);
o2 : out unsigned(0 downto 0);
o3 : out unsigned(63 downto 0));
end component cf_fft_2048_16_30;
component cf_fft_2048_16_26 is
port (
clock_c : in std_logic;
i1 : in  unsigned(0 downto 0);
i2 : in  unsigned(0 downto 0);
i3 : in  unsigned(0 downto 0);
o1 : out unsigned(9 downto 0);
o2 : out unsigned(0 downto 0));
end component cf_fft_2048_16_26;
begin
n1 <= s29_1(9 downto 9) &
  s29_1(8 downto 8) &
  s29_1(7 downto 7) &
  s29_1(6 downto 6) &
  s29_1(5 downto 5) &
  s29_1(4 downto 4) &
  s29_1(3 downto 3) &
  s29_1(2 downto 2);
n2 <= s25_1 & s25_2;
process (clock_c) begin
  if rising_edge(clock_c) then
    if i5 = "1" then
      n3 <= "0";
    elsif i4 = "1" then
      n3 <= s29_2;
    end if;
  end if;
end process;
process (clock_c) begin
  if rising_edge(clock_c) then
    if i5 = "1" then
      n4 <= "0";
    elsif i4 = "1" then
      n4 <= n3;
    end if;
  end if;
end process;
process (clock_c) begin
  if rising_edge(clock_c) then
    if i5 = "1" then
      n5 <= "0";
    elsif i4 = "1" then
      n5 <= n4;
    end if;
  end if;
end process;
process (clock_c) begin
  if rising_edge(clock_c) then
    if i5 = "1" then
      n6 <= "0";
    elsif i4 = "1" then
      n6 <= n5;
    end if;
  end if;
end process;
n7 <= s29_1(9 downto 9) &
  s29_1(8 downto 8) &
  s29_1(7 downto 7) &
  s29_1(6 downto 6) &
  s29_1(5 downto 5) &
  s29_1(4 downto 4) &
  s29_1(3 downto 3) &
  s29_1(2 downto 2) &
  s29_1(1 downto 1);
process (clock_c) begin
  if rising_edge(clock_c) then
    if i5 = "1" then
      n8 <= "000000000";
    elsif i4 = "1" then
      n8 <= n7;
    end if;
  end if;
end process;
process (clock_c) begin
  if rising_edge(clock_c) then
    if i5 = "1" then
      n9 <= "000000000";
    elsif i4 = "1" then
      n9 <= n8;
    end if;
  end if;
end process;
process (clock_c) begin
  if rising_edge(clock_c) then
    if i5 = "1" then
      n10 <= "000000000";
    elsif i4 = "1" then
      n10 <= n9;
    end if;
  end if;
end process;
process (clock_c) begin
  if rising_edge(clock_c) then
    if i5 = "1" then
      n11 <= "000000000";
    elsif i4 = "1" then
      n11 <= n10;
    end if;
  end if;
end process;
n12 <= s29_1(0 downto 0);
process (clock_c) begin
  if rising_edge(clock_c) then
    if i5 = "1" then
      n13 <= "0";
    elsif i4 = "1" then
      n13 <= n12;
    end if;
  end if;
end process;
process (clock_c) begin
  if rising_edge(clock_c) then
    if i5 = "1" then
      n14 <= "0";
    elsif i4 = "1" then
      n14 <= n13;
    end if;
  end if;
end process;
process (clock_c) begin
  if rising_edge(clock_c) then
    if i5 = "1" then
      n15 <= "0";
    elsif i4 = "1" then
      n15 <= n14;
    end if;
  end if;
end process;
process (clock_c) begin
  if rising_edge(clock_c) then
    if i5 = "1" then
      n16 <= "0";
    elsif i4 = "1" then
      n16 <= n15;
    end if;
  end if;
end process;
n17 <= not n16;
n18 <= s28_2 & s28_1;
n19 <= s28_3(63 downto 63) &
  s28_3(62 downto 62) &
  s28_3(61 downto 61) &
  s28_3(60 downto 60) &
  s28_3(59 downto 59) &
  s28_3(58 downto 58) &
  s28_3(57 downto 57) &
  s28_3(56 downto 56) &
  s28_3(55 downto 55) &
  s28_3(54 downto 54) &
  s28_3(53 downto 53) &
  s28_3(52 downto 52) &
  s28_3(51 downto 51) &
  s28_3(50 downto 50) &
  s28_3(49 downto 49) &
  s28_3(48 downto 48) &
  s28_3(47 downto 47) &
  s28_3(46 downto 46) &
  s28_3(45 downto 45) &
  s28_3(44 downto 44) &
  s28_3(43 downto 43) &
  s28_3(42 downto 42) &
  s28_3(41 downto 41) &
  s28_3(40 downto 40) &
  s28_3(39 downto 39) &
  s28_3(38 downto 38) &
  s28_3(37 downto 37) &
  s28_3(36 downto 36) &
  s28_3(35 downto 35) &
  s28_3(34 downto 34) &
  s28_3(33 downto 33) &
  s28_3(32 downto 32);
n20 <= s28_3(31 downto 31) &
  s28_3(30 downto 30) &
  s28_3(29 downto 29) &
  s28_3(28 downto 28) &
  s28_3(27 downto 27) &
  s28_3(26 downto 26) &
  s28_3(25 downto 25) &
  s28_3(24 downto 24) &
  s28_3(23 downto 23) &
  s28_3(22 downto 22) &
  s28_3(21 downto 21) &
  s28_3(20 downto 20) &
  s28_3(19 downto 19) &
  s28_3(18 downto 18) &
  s28_3(17 downto 17) &
  s28_3(16 downto 16) &
  s28_3(15 downto 15) &
  s28_3(14 downto 14) &
  s28_3(13 downto 13) &
  s28_3(12 downto 12) &
  s28_3(11 downto 11) &
  s28_3(10 downto 10) &
  s28_3(9 downto 9) &
  s28_3(8 downto 8) &
  s28_3(7 downto 7) &
  s28_3(6 downto 6) &
  s28_3(5 downto 5) &
  s28_3(4 downto 4) &
  s28_3(3 downto 3) &
  s28_3(2 downto 2) &
  s28_3(1 downto 1) &
  s28_3(0 downto 0);
n21 <= s27_1(63 downto 63) &
  s27_1(62 downto 62) &
  s27_1(61 downto 61) &
  s27_1(60 downto 60) &
  s27_1(59 downto 59) &
  s27_1(58 downto 58) &
  s27_1(57 downto 57) &
  s27_1(56 downto 56) &
  s27_1(55 downto 55) &
  s27_1(54 downto 54) &
  s27_1(53 downto 53) &
  s27_1(52 downto 52) &
  s27_1(51 downto 51) &
  s27_1(50 downto 50) &
  s27_1(49 downto 49) &
  s27_1(48 downto 48) &
  s27_1(47 downto 47) &
  s27_1(46 downto 46) &
  s27_1(45 downto 45) &
  s27_1(44 downto 44) &
  s27_1(43 downto 43) &
  s27_1(42 downto 42) &
  s27_1(41 downto 41) &
  s27_1(40 downto 40) &
  s27_1(39 downto 39) &
  s27_1(38 downto 38) &
  s27_1(37 downto 37) &
  s27_1(36 downto 36) &
  s27_1(35 downto 35) &
  s27_1(34 downto 34) &
  s27_1(33 downto 33) &
  s27_1(32 downto 32);
n22 <= s27_1(31 downto 31) &
  s27_1(30 downto 30) &
  s27_1(29 downto 29) &
  s27_1(28 downto 28) &
  s27_1(27 downto 27) &
  s27_1(26 downto 26) &
  s27_1(25 downto 25) &
  s27_1(24 downto 24) &
  s27_1(23 downto 23) &
  s27_1(22 downto 22) &
  s27_1(21 downto 21) &
  s27_1(20 downto 20) &
  s27_1(19 downto 19) &
  s27_1(18 downto 18) &
  s27_1(17 downto 17) &
  s27_1(16 downto 16) &
  s27_1(15 downto 15) &
  s27_1(14 downto 14) &
  s27_1(13 downto 13) &
  s27_1(12 downto 12) &
  s27_1(11 downto 11) &
  s27_1(10 downto 10) &
  s27_1(9 downto 9) &
  s27_1(8 downto 8) &
  s27_1(7 downto 7) &
  s27_1(6 downto 6) &
  s27_1(5 downto 5) &
  s27_1(4 downto 4) &
  s27_1(3 downto 3) &
  s27_1(2 downto 2) &
  s27_1(1 downto 1) &
  s27_1(0 downto 0);
n23 <= n20 when s26_1 = "1" else n19;
n24 <= n22 when s26_1 = "1" else n21;
s25 : cf_fft_2048_16_20 port map (clock_c, i2, i3, n1, i4, i5, s25_1, s25_2);
s26 : cf_fft_2048_16_35 port map (clock_c, n18, i4, i5, s26_1);
s27 : cf_fft_2048_16_31 port map (clock_c, n2, n6, n11, n16, i4, i5, s27_1);
s28 : cf_fft_2048_16_30 port map (clock_c, n2, n6, n11, n17, i4, i5, s28_1, s28_2, s28_3);
s29 : cf_fft_2048_16_26 port map (clock_c, i1, i4, i5, s29_1, s29_2);
o3 <= n24;
o2 <= n23;
o1 <= s28_1;
end architecture rtl;

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
entity cf_fft_2048_16_18 is
port (
clock_c : in std_logic;
i1 : in  unsigned(31 downto 0);
i2 : in  unsigned(31 downto 0);
i3 : in  unsigned(6 downto 0);
i4 : in  unsigned(0 downto 0);
i5 : in  unsigned(0 downto 0);
o1 : out unsigned(31 downto 0);
o2 : out unsigned(31 downto 0));
end entity cf_fft_2048_16_18;
architecture rtl of cf_fft_2048_16_18 is
signal n1 : unsigned(31 downto 0) := "00000000000000000000000000000000";
signal n2 : unsigned(15 downto 0);
signal n3 : unsigned(15 downto 0);
signal n4 : unsigned(31 downto 0) := "00000000000000000000000000000000";
signal n5 : unsigned(15 downto 0);
signal n6 : unsigned(15 downto 0);
signal n7 : unsigned(15 downto 0) := "0000000000000000";
signal n8 : unsigned(15 downto 0) := "0000000000000000";
signal n9 : unsigned(15 downto 0) := "0000000000000000";
signal n10 : unsigned(15 downto 0) := "0000000000000000";
signal n11 : unsigned(31 downto 0) := "00000000000000000000000000000000";
signal n12 : unsigned(15 downto 0);
signal n13 : unsigned(15 downto 0);
signal n14 : unsigned(31 downto 0);
signal n15 : unsigned(15 downto 0);
signal n16 : unsigned(15 downto 0) := "0000000000000000";
signal n17 : unsigned(31 downto 0);
signal n18 : unsigned(15 downto 0);
signal n19 : unsigned(15 downto 0) := "0000000000000000";
signal n20 : unsigned(15 downto 0);
signal n21 : unsigned(15 downto 0) := "0000000000000000";
signal n22 : unsigned(31 downto 0);
signal n23 : unsigned(15 downto 0);
signal n24 : unsigned(15 downto 0) := "0000000000000000";
signal n25 : unsigned(31 downto 0);
signal n26 : unsigned(15 downto 0);
signal n27 : unsigned(15 downto 0) := "0000000000000000";
signal n28 : unsigned(15 downto 0);
signal n29 : unsigned(15 downto 0) := "0000000000000000";
signal n30 : unsigned(15 downto 0);
signal n31 : unsigned(15 downto 0);
signal n32 : unsigned(31 downto 0);
signal n33 : unsigned(31 downto 0) := "00000000000000000000000000000000";
signal n34 : unsigned(15 downto 0);
signal n35 : unsigned(15 downto 0);
signal n36 : unsigned(31 downto 0);
signal n37 : unsigned(31 downto 0) := "00000000000000000000000000000000";
begin
process (clock_c) begin
  if rising_edge(clock_c) then
    if i5 = "1" then
      n1 <= "00000000000000000000000000000000";
    elsif i4 = "1" then
      n1 <= i1;
    end if;
  end if;
end process;
n2 <= n1(31 downto 31) &
  n1(30 downto 30) &
  n1(29 downto 29) &
  n1(28 downto 28) &
  n1(27 downto 27) &
  n1(26 downto 26) &
  n1(25 downto 25) &
  n1(24 downto 24) &
  n1(23 downto 23) &
  n1(22 downto 22) &
  n1(21 downto 21) &
  n1(20 downto 20) &
  n1(19 downto 19) &
  n1(18 downto 18) &
  n1(17 downto 17) &
  n1(16 downto 16);
n3 <= n1(15 downto 15) &
  n1(14 downto 14) &
  n1(13 downto 13) &
  n1(12 downto 12) &
  n1(11 downto 11) &
  n1(10 downto 10) &
  n1(9 downto 9) &
  n1(8 downto 8) &
  n1(7 downto 7) &
  n1(6 downto 6) &
  n1(5 downto 5) &
  n1(4 downto 4) &
  n1(3 downto 3) &
  n1(2 downto 2) &
  n1(1 downto 1) &
  n1(0 downto 0);
process (clock_c) begin
  if rising_edge(clock_c) then
    if i5 = "1" then
      n4 <= "00000000000000000000000000000000";
    elsif i4 = "1" then
      n4 <= i2;
    end if;
  end if;
end process;
n5 <= n4(31 downto 31) &
  n4(30 downto 30) &
  n4(29 downto 29) &
  n4(28 downto 28) &
  n4(27 downto 27) &
  n4(26 downto 26) &
  n4(25 downto 25) &
  n4(24 downto 24) &
  n4(23 downto 23) &
  n4(22 downto 22) &
  n4(21 downto 21) &
  n4(20 downto 20) &
  n4(19 downto 19) &
  n4(18 downto 18) &
  n4(17 downto 17) &
  n4(16 downto 16);
n6 <= n4(15 downto 15) &
  n4(14 downto 14) &
  n4(13 downto 13) &
  n4(12 downto 12) &
  n4(11 downto 11) &
  n4(10 downto 10) &
  n4(9 downto 9) &
  n4(8 downto 8) &
  n4(7 downto 7) &
  n4(6 downto 6) &
  n4(5 downto 5) &
  n4(4 downto 4) &
  n4(3 downto 3) &
  n4(2 downto 2) &
  n4(1 downto 1) &
  n4(0 downto 0);
process (clock_c) begin
  if rising_edge(clock_c) then
    if i5 = "1" then
      n7 <= "0000000000000000";
    elsif i4 = "1" then
      n7 <= n2;
    end if;
  end if;
end process;
process (clock_c) begin
  if rising_edge(clock_c) then
    if i5 = "1" then
      n8 <= "0000000000000000";
    elsif i4 = "1" then
      n8 <= n7;
    end if;
  end if;
end process;
process (clock_c) begin
  if rising_edge(clock_c) then
    if i5 = "1" then
      n9 <= "0000000000000000";
    elsif i4 = "1" then
      n9 <= n3;
    end if;
  end if;
end process;
process (clock_c) begin
  if rising_edge(clock_c) then
    if i5 = "1" then
      n10 <= "0000000000000000";
    elsif i4 = "1" then
      n10 <= n9;
    end if;
  end if;
end process;
process (clock_c) begin
  if rising_edge(clock_c) then 
    if i4 = "1" then
      case i3 is
        when "0000000" => n11 <= "01111111111111110000000000000000";
        when "0000001" => n11 <= "01111111111101101111110011011011";
        when "0000010" => n11 <= "01111111110110001111100110111000";
        when "0000011" => n11 <= "01111111101001111111011010010101";
        when "0000100" => n11 <= "01111111011000101111001101110100";
        when "0000101" => n11 <= "01111111000010011111000001010100";
        when "0000110" => n11 <= "01111110100111011110110100110111";
        when "0000111" => n11 <= "01111110000111011110101000011101";
        when "0001000" => n11 <= "01111101100010101110011100000111";
        when "0001001" => n11 <= "01111100111000111110001111110100";
        when "0001010" => n11 <= "01111100001010011110000011100110";
        when "0001011" => n11 <= "01111011010111011101110111011100";
        when "0001100" => n11 <= "01111010011111011101101011010111";
        when "0001101" => n11 <= "01111001100010101101011111011001";
        when "0001110" => n11 <= "01111000100001001101010011100000";
        when "0001111" => n11 <= "01110111011011001101000111101110";
        when "0010000" => n11 <= "01110110010000011100111100000100";
        when "0010001" => n11 <= "01110101000001001100110000100001";
        when "0010010" => n11 <= "01110011101101011100100101000101";
        when "0010011" => n11 <= "01110010010101011100011001110011";
        when "0010100" => n11 <= "01110000111000101100001110101001";
        when "0010101" => n11 <= "01101111010111111100000011101000";
        when "0010110" => n11 <= "01101101110010101011111000110001";
        when "0010111" => n11 <= "01101100001001001011101110000101";
        when "0011000" => n11 <= "01101010011011011011100011100011";
        when "0011001" => n11 <= "01101000101001101011011001001011";
        when "0011010" => n11 <= "01100110110011111011001111000000";
        when "0011011" => n11 <= "01100100111010001011000101000000";
        when "0011100" => n11 <= "01100010111100101010111011001100";
        when "0011101" => n11 <= "01100000111011001010110001100100";
        when "0011110" => n11 <= "01011110110101111010101000001010";
        when "0011111" => n11 <= "01011100101101001010011110111101";
        when "0100000" => n11 <= "01011010100000101010010101111101";
        when "0100001" => n11 <= "01011000010000101010001101001011";
        when "0100010" => n11 <= "01010101111101011010000100101000";
        when "0100011" => n11 <= "01010011100110111001111100010011";
        when "0100100" => n11 <= "01010001001100111001110100001101";
        when "0100101" => n11 <= "01001110101111111001101100010111";
        when "0100110" => n11 <= "01001100001111111001100100110000";
        when "0100111" => n11 <= "01001001101101001001011101011001";
        when "0101000" => n11 <= "01000111000111001001010110010010";
        when "0101001" => n11 <= "01000100011110101001001111011011";
        when "0101010" => n11 <= "01000001110011101001001000110101";
        when "0101011" => n11 <= "00111111000101111001000010100000";
        when "0101100" => n11 <= "00111100010101101000111100011101";
        when "0101101" => n11 <= "00111001100011001000110110101010";
        when "0101110" => n11 <= "00110110101110101000110001001010";
        when "0101111" => n11 <= "00110011110111101000101011111011";
        when "0110000" => n11 <= "00110000111110111000100110111110";
        when "0110001" => n11 <= "00101110000100011000100010010011";
        when "0110010" => n11 <= "00101011000111111000011101111011";
        when "0110011" => n11 <= "00101000001001101000011001110101";
        when "0110100" => n11 <= "00100101001010001000010110000010";
        when "0110101" => n11 <= "00100010001000111000010010100010";
        when "0110110" => n11 <= "00011111000110011000001111010110";
        when "0110111" => n11 <= "00011100000010111000001100011100";
        when "0111000" => n11 <= "00011000111110001000001001110101";
        when "0111001" => n11 <= "00010101111000101000000111100010";
        when "0111010" => n11 <= "00010010110010001000000101100010";
        when "0111011" => n11 <= "00001111101010111000000011110110";
        when "0111100" => n11 <= "00001100100010111000000010011101";
        when "0111101" => n11 <= "00001001011010101000000001011000";
        when "0111110" => n11 <= "00000110010001111000000000100111";
        when "0111111" => n11 <= "00000011001001001000000000001001";
        when "1000000" => n11 <= "00000000000000001000000000000000";
        when "1000001" => n11 <= "11111100110110111000000000001001";
        when "1000010" => n11 <= "11111001101110001000000000100111";
        when "1000011" => n11 <= "11110110100101011000000001011000";
        when "1000100" => n11 <= "11110011011101001000000010011101";
        when "1000101" => n11 <= "11110000010101001000000011110110";
        when "1000110" => n11 <= "11101101001101111000000101100010";
        when "1000111" => n11 <= "11101010000111011000000111100010";
        when "1001000" => n11 <= "11100111000001111000001001110101";
        when "1001001" => n11 <= "11100011111101001000001100011100";
        when "1001010" => n11 <= "11100000111001101000001111010110";
        when "1001011" => n11 <= "11011101110111001000010010100010";
        when "1001100" => n11 <= "11011010110101111000010110000010";
        when "1001101" => n11 <= "11010111110110011000011001110101";
        when "1001110" => n11 <= "11010100111000001000011101111011";
        when "1001111" => n11 <= "11010001111011101000100010010011";
        when "1010000" => n11 <= "11001111000001001000100110111110";
        when "1010001" => n11 <= "11001100001000011000101011111011";
        when "1010010" => n11 <= "11001001010001011000110001001010";
        when "1010011" => n11 <= "11000110011100111000110110101010";
        when "1010100" => n11 <= "11000011101010011000111100011101";
        when "1010101" => n11 <= "11000000111010001001000010100000";
        when "1010110" => n11 <= "10111110001100011001001000110101";
        when "1010111" => n11 <= "10111011100001011001001111011011";
        when "1011000" => n11 <= "10111000111000111001010110010010";
        when "1011001" => n11 <= "10110110010010111001011101011001";
        when "1011010" => n11 <= "10110011110000001001100100110000";
        when "1011011" => n11 <= "10110001010000001001101100010111";
        when "1011100" => n11 <= "10101110110011001001110100001101";
        when "1011101" => n11 <= "10101100011001001001111100010011";
        when "1011110" => n11 <= "10101010000010101010000100101000";
        when "1011111" => n11 <= "10100111101111011010001101001011";
        when "1100000" => n11 <= "10100101011111011010010101111101";
        when "1100001" => n11 <= "10100011010010111010011110111101";
        when "1100010" => n11 <= "10100001001010001010101000001010";
        when "1100011" => n11 <= "10011111000100111010110001100100";
        when "1100100" => n11 <= "10011101000011011010111011001100";
        when "1100101" => n11 <= "10011011000101111011000101000000";
        when "1100110" => n11 <= "10011001001100001011001111000000";
        when "1100111" => n11 <= "10010111010110011011011001001011";
        when "1101000" => n11 <= "10010101100100101011100011100011";
        when "1101001" => n11 <= "10010011110110111011101110000101";
        when "1101010" => n11 <= "10010010001101011011111000110001";
        when "1101011" => n11 <= "10010000101000001100000011101000";
        when "1101100" => n11 <= "10001111000111011100001110101001";
        when "1101101" => n11 <= "10001101101010101100011001110011";
        when "1101110" => n11 <= "10001100010010101100100101000101";
        when "1101111" => n11 <= "10001010111110111100110000100001";
        when "1110000" => n11 <= "10001001101111101100111100000100";
        when "1110001" => n11 <= "10001000100100111101000111101110";
        when "1110010" => n11 <= "10000111011110111101010011100000";
        when "1110011" => n11 <= "10000110011101011101011111011001";
        when "1110100" => n11 <= "10000101100000101101101011010111";
        when "1110101" => n11 <= "10000100101000101101110111011100";
        when "1110110" => n11 <= "10000011110101101110000011100110";
        when "1110111" => n11 <= "10000011000111001110001111110100";
        when "1111000" => n11 <= "10000010011101011110011100000111";
        when "1111001" => n11 <= "10000001111000101110101000011101";
        when "1111010" => n11 <= "10000001011000101110110100110111";
        when "1111011" => n11 <= "10000000111101101111000001010100";
        when "1111100" => n11 <= "10000000100111011111001101110100";
        when "1111101" => n11 <= "10000000010110001111011010010101";
        when "1111110" => n11 <= "10000000001001111111100110111000";
        when "1111111" => n11 <= "10000000000010011111110011011011";
        when others => n11 <= "XXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX";
      end case;
    end if;
  end if;
end process;
n12 <= n11(31 downto 31) &
  n11(30 downto 30) &
  n11(29 downto 29) &
  n11(28 downto 28) &
  n11(27 downto 27) &
  n11(26 downto 26) &
  n11(25 downto 25) &
  n11(24 downto 24) &
  n11(23 downto 23) &
  n11(22 downto 22) &
  n11(21 downto 21) &
  n11(20 downto 20) &
  n11(19 downto 19) &
  n11(18 downto 18) &
  n11(17 downto 17) &
  n11(16 downto 16);
n13 <= n11(15 downto 15) &
  n11(14 downto 14) &
  n11(13 downto 13) &
  n11(12 downto 12) &
  n11(11 downto 11) &
  n11(10 downto 10) &
  n11(9 downto 9) &
  n11(8 downto 8) &
  n11(7 downto 7) &
  n11(6 downto 6) &
  n11(5 downto 5) &
  n11(4 downto 4) &
  n11(3 downto 3) &
  n11(2 downto 2) &
  n11(1 downto 1) &
  n11(0 downto 0);
n14 <= unsigned(signed(n5) * signed(n12));
n15 <= n14(30 downto 30) &
  n14(29 downto 29) &
  n14(28 downto 28) &
  n14(27 downto 27) &
  n14(26 downto 26) &
  n14(25 downto 25) &
  n14(24 downto 24) &
  n14(23 downto 23) &
  n14(22 downto 22) &
  n14(21 downto 21) &
  n14(20 downto 20) &
  n14(19 downto 19) &
  n14(18 downto 18) &
  n14(17 downto 17) &
  n14(16 downto 16) &
  n14(15 downto 15);
process (clock_c) begin
  if rising_edge(clock_c) then
    if i5 = "1" then
      n16 <= "0000000000000000";
    elsif i4 = "1" then
      n16 <= n15;
    end if;
  end if;
end process;
n17 <= unsigned(signed(n6) * signed(n13));
n18 <= n17(30 downto 30) &
  n17(29 downto 29) &
  n17(28 downto 28) &
  n17(27 downto 27) &
  n17(26 downto 26) &
  n17(25 downto 25) &
  n17(24 downto 24) &
  n17(23 downto 23) &
  n17(22 downto 22) &
  n17(21 downto 21) &
  n17(20 downto 20) &
  n17(19 downto 19) &
  n17(18 downto 18) &
  n17(17 downto 17) &
  n17(16 downto 16) &
  n17(15 downto 15);
process (clock_c) begin
  if rising_edge(clock_c) then
    if i5 = "1" then
      n19 <= "0000000000000000";
    elsif i4 = "1" then
      n19 <= n18;
    end if;
  end if;
end process;
n20 <= n16 - n19;
process (clock_c) begin
  if rising_edge(clock_c) then
    if i5 = "1" then
      n21 <= "0000000000000000";
    elsif i4 = "1" then
      n21 <= n20;
    end if;
  end if;
end process;
n22 <= unsigned(signed(n5) * signed(n13));
n23 <= n22(30 downto 30) &
  n22(29 downto 29) &
  n22(28 downto 28) &
  n22(27 downto 27) &
  n22(26 downto 26) &
  n22(25 downto 25) &
  n22(24 downto 24) &
  n22(23 downto 23) &
  n22(22 downto 22) &
  n22(21 downto 21) &
  n22(20 downto 20) &
  n22(19 downto 19) &
  n22(18 downto 18) &
  n22(17 downto 17) &
  n22(16 downto 16) &
  n22(15 downto 15);
process (clock_c) begin
  if rising_edge(clock_c) then
    if i5 = "1" then
      n24 <= "0000000000000000";
    elsif i4 = "1" then
      n24 <= n23;
    end if;
  end if;
end process;
n25 <= unsigned(signed(n6) * signed(n12));
n26 <= n25(30 downto 30) &
  n25(29 downto 29) &
  n25(28 downto 28) &
  n25(27 downto 27) &
  n25(26 downto 26) &
  n25(25 downto 25) &
  n25(24 downto 24) &
  n25(23 downto 23) &
  n25(22 downto 22) &
  n25(21 downto 21) &
  n25(20 downto 20) &
  n25(19 downto 19) &
  n25(18 downto 18) &
  n25(17 downto 17) &
  n25(16 downto 16) &
  n25(15 downto 15);
process (clock_c) begin
  if rising_edge(clock_c) then
    if i5 = "1" then
      n27 <= "0000000000000000";
    elsif i4 = "1" then
      n27 <= n26;
    end if;
  end if;
end process;
n28 <= n24 + n27;
process (clock_c) begin
  if rising_edge(clock_c) then
    if i5 = "1" then
      n29 <= "0000000000000000";
    elsif i4 = "1" then
      n29 <= n28;
    end if;
  end if;
end process;
n30 <= n8 + n21;
n31 <= n10 + n29;
n32 <= n30 & n31;
process (clock_c) begin
  if rising_edge(clock_c) then
    if i5 = "1" then
      n33 <= "00000000000000000000000000000000";
    elsif i4 = "1" then
      n33 <= n32;
    end if;
  end if;
end process;
n34 <= n8 - n21;
n35 <= n10 - n29;
n36 <= n34 & n35;
process (clock_c) begin
  if rising_edge(clock_c) then
    if i5 = "1" then
      n37 <= "00000000000000000000000000000000";
    elsif i4 = "1" then
      n37 <= n36;
    end if;
  end if;
end process;
o2 <= n37;
o1 <= n33;
end architecture rtl;

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
entity cf_fft_2048_16_17 is
port (
clock_c : in std_logic;
i1 : in  unsigned(0 downto 0);
i2 : in  unsigned(31 downto 0);
i3 : in  unsigned(31 downto 0);
i4 : in  unsigned(0 downto 0);
i5 : in  unsigned(0 downto 0);
o1 : out unsigned(0 downto 0);
o2 : out unsigned(31 downto 0);
o3 : out unsigned(31 downto 0));
end entity cf_fft_2048_16_17;
architecture rtl of cf_fft_2048_16_17 is
signal n1 : unsigned(6 downto 0);
signal n2 : unsigned(63 downto 0);
signal n3 : unsigned(0 downto 0) := "0";
signal n4 : unsigned(0 downto 0) := "0";
signal n5 : unsigned(0 downto 0) := "0";
signal n6 : unsigned(0 downto 0) := "0";
signal n7 : unsigned(8 downto 0);
signal n8 : unsigned(8 downto 0) := "000000000";
signal n9 : unsigned(8 downto 0) := "000000000";
signal n10 : unsigned(8 downto 0) := "000000000";
signal n11 : unsigned(8 downto 0) := "000000000";
signal n12 : unsigned(0 downto 0);
signal n13 : unsigned(0 downto 0) := "0";
signal n14 : unsigned(0 downto 0) := "0";
signal n15 : unsigned(0 downto 0) := "0";
signal n16 : unsigned(0 downto 0) := "0";
signal n17 : unsigned(0 downto 0);
signal n18 : unsigned(1 downto 0);
signal n19 : unsigned(31 downto 0);
signal n20 : unsigned(31 downto 0);
signal n21 : unsigned(31 downto 0);
signal n22 : unsigned(31 downto 0);
signal n23 : unsigned(31 downto 0);
signal n24 : unsigned(31 downto 0);
signal s25_1 : unsigned(31 downto 0);
signal s25_2 : unsigned(31 downto 0);
signal s26_1 : unsigned(0 downto 0);
signal s27_1 : unsigned(9 downto 0);
signal s27_2 : unsigned(0 downto 0);
signal s28_1 : unsigned(63 downto 0);
signal s29_1 : unsigned(0 downto 0);
signal s29_2 : unsigned(0 downto 0);
signal s29_3 : unsigned(63 downto 0);
component cf_fft_2048_16_18 is
port (
clock_c : in std_logic;
i1 : in  unsigned(31 downto 0);
i2 : in  unsigned(31 downto 0);
i3 : in  unsigned(6 downto 0);
i4 : in  unsigned(0 downto 0);
i5 : in  unsigned(0 downto 0);
o1 : out unsigned(31 downto 0);
o2 : out unsigned(31 downto 0));
end component cf_fft_2048_16_18;
component cf_fft_2048_16_35 is
port (
clock_c : in std_logic;
i1 : in  unsigned(1 downto 0);
i2 : in  unsigned(0 downto 0);
i3 : in  unsigned(0 downto 0);
o1 : out unsigned(0 downto 0));
end component cf_fft_2048_16_35;
component cf_fft_2048_16_26 is
port (
clock_c : in std_logic;
i1 : in  unsigned(0 downto 0);
i2 : in  unsigned(0 downto 0);
i3 : in  unsigned(0 downto 0);
o1 : out unsigned(9 downto 0);
o2 : out unsigned(0 downto 0));
end component cf_fft_2048_16_26;
component cf_fft_2048_16_31 is
port (
clock_c : in std_logic;
i1 : in  unsigned(63 downto 0);
i2 : in  unsigned(0 downto 0);
i3 : in  unsigned(8 downto 0);
i4 : in  unsigned(0 downto 0);
i5 : in  unsigned(0 downto 0);
i6 : in  unsigned(0 downto 0);
o1 : out unsigned(63 downto 0));
end component cf_fft_2048_16_31;
component cf_fft_2048_16_30 is
port (
clock_c : in std_logic;
i1 : in  unsigned(63 downto 0);
i2 : in  unsigned(0 downto 0);
i3 : in  unsigned(8 downto 0);
i4 : in  unsigned(0 downto 0);
i5 : in  unsigned(0 downto 0);
i6 : in  unsigned(0 downto 0);
o1 : out unsigned(0 downto 0);
o2 : out unsigned(0 downto 0);
o3 : out unsigned(63 downto 0));
end component cf_fft_2048_16_30;
begin
n1 <= s27_1(9 downto 9) &
  s27_1(8 downto 8) &
  s27_1(7 downto 7) &
  s27_1(6 downto 6) &
  s27_1(5 downto 5) &
  s27_1(4 downto 4) &
  s27_1(3 downto 3);
n2 <= s25_1 & s25_2;
process (clock_c) begin
  if rising_edge(clock_c) then
    if i5 = "1" then
      n3 <= "0";
    elsif i4 = "1" then
      n3 <= s27_2;
    end if;
  end if;
end process;
process (clock_c) begin
  if rising_edge(clock_c) then
    if i5 = "1" then
      n4 <= "0";
    elsif i4 = "1" then
      n4 <= n3;
    end if;
  end if;
end process;
process (clock_c) begin
  if rising_edge(clock_c) then
    if i5 = "1" then
      n5 <= "0";
    elsif i4 = "1" then
      n5 <= n4;
    end if;
  end if;
end process;
process (clock_c) begin
  if rising_edge(clock_c) then
    if i5 = "1" then
      n6 <= "0";
    elsif i4 = "1" then
      n6 <= n5;
    end if;
  end if;
end process;
n7 <= s27_1(9 downto 9) &
  s27_1(8 downto 8) &
  s27_1(7 downto 7) &
  s27_1(6 downto 6) &
  s27_1(5 downto 5) &
  s27_1(4 downto 4) &
  s27_1(3 downto 3) &
  s27_1(2 downto 2) &
  s27_1(1 downto 1);
process (clock_c) begin
  if rising_edge(clock_c) then
    if i5 = "1" then
      n8 <= "000000000";
    elsif i4 = "1" then
      n8 <= n7;
    end if;
  end if;
end process;
process (clock_c) begin
  if rising_edge(clock_c) then
    if i5 = "1" then
      n9 <= "000000000";
    elsif i4 = "1" then
      n9 <= n8;
    end if;
  end if;
end process;
process (clock_c) begin
  if rising_edge(clock_c) then
    if i5 = "1" then
      n10 <= "000000000";
    elsif i4 = "1" then
      n10 <= n9;
    end if;
  end if;
end process;
process (clock_c) begin
  if rising_edge(clock_c) then
    if i5 = "1" then
      n11 <= "000000000";
    elsif i4 = "1" then
      n11 <= n10;
    end if;
  end if;
end process;
n12 <= s27_1(0 downto 0);
process (clock_c) begin
  if rising_edge(clock_c) then
    if i5 = "1" then
      n13 <= "0";
    elsif i4 = "1" then
      n13 <= n12;
    end if;
  end if;
end process;
process (clock_c) begin
  if rising_edge(clock_c) then
    if i5 = "1" then
      n14 <= "0";
    elsif i4 = "1" then
      n14 <= n13;
    end if;
  end if;
end process;
process (clock_c) begin
  if rising_edge(clock_c) then
    if i5 = "1" then
      n15 <= "0";
    elsif i4 = "1" then
      n15 <= n14;
    end if;
  end if;
end process;
process (clock_c) begin
  if rising_edge(clock_c) then
    if i5 = "1" then
      n16 <= "0";
    elsif i4 = "1" then
      n16 <= n15;
    end if;
  end if;
end process;
n17 <= not n16;
n18 <= s29_2 & s29_1;
n19 <= s29_3(63 downto 63) &
  s29_3(62 downto 62) &
  s29_3(61 downto 61) &
  s29_3(60 downto 60) &
  s29_3(59 downto 59) &
  s29_3(58 downto 58) &
  s29_3(57 downto 57) &
  s29_3(56 downto 56) &
  s29_3(55 downto 55) &
  s29_3(54 downto 54) &
  s29_3(53 downto 53) &
  s29_3(52 downto 52) &
  s29_3(51 downto 51) &
  s29_3(50 downto 50) &
  s29_3(49 downto 49) &
  s29_3(48 downto 48) &
  s29_3(47 downto 47) &
  s29_3(46 downto 46) &
  s29_3(45 downto 45) &
  s29_3(44 downto 44) &
  s29_3(43 downto 43) &
  s29_3(42 downto 42) &
  s29_3(41 downto 41) &
  s29_3(40 downto 40) &
  s29_3(39 downto 39) &
  s29_3(38 downto 38) &
  s29_3(37 downto 37) &
  s29_3(36 downto 36) &
  s29_3(35 downto 35) &
  s29_3(34 downto 34) &
  s29_3(33 downto 33) &
  s29_3(32 downto 32);
n20 <= s29_3(31 downto 31) &
  s29_3(30 downto 30) &
  s29_3(29 downto 29) &
  s29_3(28 downto 28) &
  s29_3(27 downto 27) &
  s29_3(26 downto 26) &
  s29_3(25 downto 25) &
  s29_3(24 downto 24) &
  s29_3(23 downto 23) &
  s29_3(22 downto 22) &
  s29_3(21 downto 21) &
  s29_3(20 downto 20) &
  s29_3(19 downto 19) &
  s29_3(18 downto 18) &
  s29_3(17 downto 17) &
  s29_3(16 downto 16) &
  s29_3(15 downto 15) &
  s29_3(14 downto 14) &
  s29_3(13 downto 13) &
  s29_3(12 downto 12) &
  s29_3(11 downto 11) &
  s29_3(10 downto 10) &
  s29_3(9 downto 9) &
  s29_3(8 downto 8) &
  s29_3(7 downto 7) &
  s29_3(6 downto 6) &
  s29_3(5 downto 5) &
  s29_3(4 downto 4) &
  s29_3(3 downto 3) &
  s29_3(2 downto 2) &
  s29_3(1 downto 1) &
  s29_3(0 downto 0);
n21 <= s28_1(63 downto 63) &
  s28_1(62 downto 62) &
  s28_1(61 downto 61) &
  s28_1(60 downto 60) &
  s28_1(59 downto 59) &
  s28_1(58 downto 58) &
  s28_1(57 downto 57) &
  s28_1(56 downto 56) &
  s28_1(55 downto 55) &
  s28_1(54 downto 54) &
  s28_1(53 downto 53) &
  s28_1(52 downto 52) &
  s28_1(51 downto 51) &
  s28_1(50 downto 50) &
  s28_1(49 downto 49) &
  s28_1(48 downto 48) &
  s28_1(47 downto 47) &
  s28_1(46 downto 46) &
  s28_1(45 downto 45) &
  s28_1(44 downto 44) &
  s28_1(43 downto 43) &
  s28_1(42 downto 42) &
  s28_1(41 downto 41) &
  s28_1(40 downto 40) &
  s28_1(39 downto 39) &
  s28_1(38 downto 38) &
  s28_1(37 downto 37) &
  s28_1(36 downto 36) &
  s28_1(35 downto 35) &
  s28_1(34 downto 34) &
  s28_1(33 downto 33) &
  s28_1(32 downto 32);
n22 <= s28_1(31 downto 31) &
  s28_1(30 downto 30) &
  s28_1(29 downto 29) &
  s28_1(28 downto 28) &
  s28_1(27 downto 27) &
  s28_1(26 downto 26) &
  s28_1(25 downto 25) &
  s28_1(24 downto 24) &
  s28_1(23 downto 23) &
  s28_1(22 downto 22) &
  s28_1(21 downto 21) &
  s28_1(20 downto 20) &
  s28_1(19 downto 19) &
  s28_1(18 downto 18) &
  s28_1(17 downto 17) &
  s28_1(16 downto 16) &
  s28_1(15 downto 15) &
  s28_1(14 downto 14) &
  s28_1(13 downto 13) &
  s28_1(12 downto 12) &
  s28_1(11 downto 11) &
  s28_1(10 downto 10) &
  s28_1(9 downto 9) &
  s28_1(8 downto 8) &
  s28_1(7 downto 7) &
  s28_1(6 downto 6) &
  s28_1(5 downto 5) &
  s28_1(4 downto 4) &
  s28_1(3 downto 3) &
  s28_1(2 downto 2) &
  s28_1(1 downto 1) &
  s28_1(0 downto 0);
n23 <= n20 when s26_1 = "1" else n19;
n24 <= n22 when s26_1 = "1" else n21;
s25 : cf_fft_2048_16_18 port map (clock_c, i2, i3, n1, i4, i5, s25_1, s25_2);
s26 : cf_fft_2048_16_35 port map (clock_c, n18, i4, i5, s26_1);
s27 : cf_fft_2048_16_26 port map (clock_c, i1, i4, i5, s27_1, s27_2);
s28 : cf_fft_2048_16_31 port map (clock_c, n2, n6, n11, n16, i4, i5, s28_1);
s29 : cf_fft_2048_16_30 port map (clock_c, n2, n6, n11, n17, i4, i5, s29_1, s29_2, s29_3);
o3 <= n24;
o2 <= n23;
o1 <= s29_1;
end architecture rtl;

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
entity cf_fft_2048_16_16 is
port (
clock_c : in std_logic;
i1 : in  unsigned(31 downto 0);
i2 : in  unsigned(31 downto 0);
i3 : in  unsigned(5 downto 0);
i4 : in  unsigned(0 downto 0);
i5 : in  unsigned(0 downto 0);
o1 : out unsigned(31 downto 0);
o2 : out unsigned(31 downto 0));
end entity cf_fft_2048_16_16;
architecture rtl of cf_fft_2048_16_16 is
signal n1 : unsigned(31 downto 0) := "00000000000000000000000000000000";
signal n2 : unsigned(15 downto 0);
signal n3 : unsigned(15 downto 0);
signal n4 : unsigned(31 downto 0) := "00000000000000000000000000000000";
signal n5 : unsigned(15 downto 0);
signal n6 : unsigned(15 downto 0);
signal n7 : unsigned(15 downto 0) := "0000000000000000";
signal n8 : unsigned(15 downto 0) := "0000000000000000";
signal n9 : unsigned(15 downto 0) := "0000000000000000";
signal n10 : unsigned(15 downto 0) := "0000000000000000";
signal n11 : unsigned(31 downto 0) := "00000000000000000000000000000000";
signal n12 : unsigned(15 downto 0);
signal n13 : unsigned(15 downto 0);
signal n14 : unsigned(31 downto 0);
signal n15 : unsigned(15 downto 0);
signal n16 : unsigned(15 downto 0) := "0000000000000000";
signal n17 : unsigned(31 downto 0);
signal n18 : unsigned(15 downto 0);
signal n19 : unsigned(15 downto 0) := "0000000000000000";
signal n20 : unsigned(15 downto 0);
signal n21 : unsigned(15 downto 0) := "0000000000000000";
signal n22 : unsigned(31 downto 0);
signal n23 : unsigned(15 downto 0);
signal n24 : unsigned(15 downto 0) := "0000000000000000";
signal n25 : unsigned(31 downto 0);
signal n26 : unsigned(15 downto 0);
signal n27 : unsigned(15 downto 0) := "0000000000000000";
signal n28 : unsigned(15 downto 0);
signal n29 : unsigned(15 downto 0) := "0000000000000000";
signal n30 : unsigned(15 downto 0);
signal n31 : unsigned(15 downto 0);
signal n32 : unsigned(31 downto 0);
signal n33 : unsigned(31 downto 0) := "00000000000000000000000000000000";
signal n34 : unsigned(15 downto 0);
signal n35 : unsigned(15 downto 0);
signal n36 : unsigned(31 downto 0);
signal n37 : unsigned(31 downto 0) := "00000000000000000000000000000000";
begin
process (clock_c) begin
  if rising_edge(clock_c) then
    if i5 = "1" then
      n1 <= "00000000000000000000000000000000";
    elsif i4 = "1" then
      n1 <= i1;
    end if;
  end if;
end process;
n2 <= n1(31 downto 31) &
  n1(30 downto 30) &
  n1(29 downto 29) &
  n1(28 downto 28) &
  n1(27 downto 27) &
  n1(26 downto 26) &
  n1(25 downto 25) &
  n1(24 downto 24) &
  n1(23 downto 23) &
  n1(22 downto 22) &
  n1(21 downto 21) &
  n1(20 downto 20) &
  n1(19 downto 19) &
  n1(18 downto 18) &
  n1(17 downto 17) &
  n1(16 downto 16);
n3 <= n1(15 downto 15) &
  n1(14 downto 14) &
  n1(13 downto 13) &
  n1(12 downto 12) &
  n1(11 downto 11) &
  n1(10 downto 10) &
  n1(9 downto 9) &
  n1(8 downto 8) &
  n1(7 downto 7) &
  n1(6 downto 6) &
  n1(5 downto 5) &
  n1(4 downto 4) &
  n1(3 downto 3) &
  n1(2 downto 2) &
  n1(1 downto 1) &
  n1(0 downto 0);
process (clock_c) begin
  if rising_edge(clock_c) then
    if i5 = "1" then
      n4 <= "00000000000000000000000000000000";
    elsif i4 = "1" then
      n4 <= i2;
    end if;
  end if;
end process;
n5 <= n4(31 downto 31) &
  n4(30 downto 30) &
  n4(29 downto 29) &
  n4(28 downto 28) &
  n4(27 downto 27) &
  n4(26 downto 26) &
  n4(25 downto 25) &
  n4(24 downto 24) &
  n4(23 downto 23) &
  n4(22 downto 22) &
  n4(21 downto 21) &
  n4(20 downto 20) &
  n4(19 downto 19) &
  n4(18 downto 18) &
  n4(17 downto 17) &
  n4(16 downto 16);
n6 <= n4(15 downto 15) &
  n4(14 downto 14) &
  n4(13 downto 13) &
  n4(12 downto 12) &
  n4(11 downto 11) &
  n4(10 downto 10) &
  n4(9 downto 9) &
  n4(8 downto 8) &
  n4(7 downto 7) &
  n4(6 downto 6) &
  n4(5 downto 5) &
  n4(4 downto 4) &
  n4(3 downto 3) &
  n4(2 downto 2) &
  n4(1 downto 1) &
  n4(0 downto 0);
process (clock_c) begin
  if rising_edge(clock_c) then
    if i5 = "1" then
      n7 <= "0000000000000000";
    elsif i4 = "1" then
      n7 <= n2;
    end if;
  end if;
end process;
process (clock_c) begin
  if rising_edge(clock_c) then
    if i5 = "1" then
      n8 <= "0000000000000000";
    elsif i4 = "1" then
      n8 <= n7;
    end if;
  end if;
end process;
process (clock_c) begin
  if rising_edge(clock_c) then
    if i5 = "1" then
      n9 <= "0000000000000000";
    elsif i4 = "1" then
      n9 <= n3;
    end if;
  end if;
end process;
process (clock_c) begin
  if rising_edge(clock_c) then
    if i5 = "1" then
      n10 <= "0000000000000000";
    elsif i4 = "1" then
      n10 <= n9;
    end if;
  end if;
end process;
process (clock_c) begin
  if rising_edge(clock_c) then 
    if i4 = "1" then
      case i3 is
        when "000000" => n11 <= "01111111111111110000000000000000";
        when "000001" => n11 <= "01111111110110001111100110111000";
        when "000010" => n11 <= "01111111011000101111001101110100";
        when "000011" => n11 <= "01111110100111011110110100110111";
        when "000100" => n11 <= "01111101100010101110011100000111";
        when "000101" => n11 <= "01111100001010011110000011100110";
        when "000110" => n11 <= "01111010011111011101101011010111";
        when "000111" => n11 <= "01111000100001001101010011100000";
        when "001000" => n11 <= "01110110010000011100111100000100";
        when "001001" => n11 <= "01110011101101011100100101000101";
        when "001010" => n11 <= "01110000111000101100001110101001";
        when "001011" => n11 <= "01101101110010101011111000110001";
        when "001100" => n11 <= "01101010011011011011100011100011";
        when "001101" => n11 <= "01100110110011111011001111000000";
        when "001110" => n11 <= "01100010111100101010111011001100";
        when "001111" => n11 <= "01011110110101111010101000001010";
        when "010000" => n11 <= "01011010100000101010010101111101";
        when "010001" => n11 <= "01010101111101011010000100101000";
        when "010010" => n11 <= "01010001001100111001110100001101";
        when "010011" => n11 <= "01001100001111111001100100110000";
        when "010100" => n11 <= "01000111000111001001010110010010";
        when "010101" => n11 <= "01000001110011101001001000110101";
        when "010110" => n11 <= "00111100010101101000111100011101";
        when "010111" => n11 <= "00110110101110101000110001001010";
        when "011000" => n11 <= "00110000111110111000100110111110";
        when "011001" => n11 <= "00101011000111111000011101111011";
        when "011010" => n11 <= "00100101001010001000010110000010";
        when "011011" => n11 <= "00011111000110011000001111010110";
        when "011100" => n11 <= "00011000111110001000001001110101";
        when "011101" => n11 <= "00010010110010001000000101100010";
        when "011110" => n11 <= "00001100100010111000000010011101";
        when "011111" => n11 <= "00000110010001111000000000100111";
        when "100000" => n11 <= "00000000000000001000000000000000";
        when "100001" => n11 <= "11111001101110001000000000100111";
        when "100010" => n11 <= "11110011011101001000000010011101";
        when "100011" => n11 <= "11101101001101111000000101100010";
        when "100100" => n11 <= "11100111000001111000001001110101";
        when "100101" => n11 <= "11100000111001101000001111010110";
        when "100110" => n11 <= "11011010110101111000010110000010";
        when "100111" => n11 <= "11010100111000001000011101111011";
        when "101000" => n11 <= "11001111000001001000100110111110";
        when "101001" => n11 <= "11001001010001011000110001001010";
        when "101010" => n11 <= "11000011101010011000111100011101";
        when "101011" => n11 <= "10111110001100011001001000110101";
        when "101100" => n11 <= "10111000111000111001010110010010";
        when "101101" => n11 <= "10110011110000001001100100110000";
        when "101110" => n11 <= "10101110110011001001110100001101";
        when "101111" => n11 <= "10101010000010101010000100101000";
        when "110000" => n11 <= "10100101011111011010010101111101";
        when "110001" => n11 <= "10100001001010001010101000001010";
        when "110010" => n11 <= "10011101000011011010111011001100";
        when "110011" => n11 <= "10011001001100001011001111000000";
        when "110100" => n11 <= "10010101100100101011100011100011";
        when "110101" => n11 <= "10010010001101011011111000110001";
        when "110110" => n11 <= "10001111000111011100001110101001";
        when "110111" => n11 <= "10001100010010101100100101000101";
        when "111000" => n11 <= "10001001101111101100111100000100";
        when "111001" => n11 <= "10000111011110111101010011100000";
        when "111010" => n11 <= "10000101100000101101101011010111";
        when "111011" => n11 <= "10000011110101101110000011100110";
        when "111100" => n11 <= "10000010011101011110011100000111";
        when "111101" => n11 <= "10000001011000101110110100110111";
        when "111110" => n11 <= "10000000100111011111001101110100";
        when "111111" => n11 <= "10000000001001111111100110111000";
        when others => n11 <= "XXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX";
      end case;
    end if;
  end if;
end process;
n12 <= n11(31 downto 31) &
  n11(30 downto 30) &
  n11(29 downto 29) &
  n11(28 downto 28) &
  n11(27 downto 27) &
  n11(26 downto 26) &
  n11(25 downto 25) &
  n11(24 downto 24) &
  n11(23 downto 23) &
  n11(22 downto 22) &
  n11(21 downto 21) &
  n11(20 downto 20) &
  n11(19 downto 19) &
  n11(18 downto 18) &
  n11(17 downto 17) &
  n11(16 downto 16);
n13 <= n11(15 downto 15) &
  n11(14 downto 14) &
  n11(13 downto 13) &
  n11(12 downto 12) &
  n11(11 downto 11) &
  n11(10 downto 10) &
  n11(9 downto 9) &
  n11(8 downto 8) &
  n11(7 downto 7) &
  n11(6 downto 6) &
  n11(5 downto 5) &
  n11(4 downto 4) &
  n11(3 downto 3) &
  n11(2 downto 2) &
  n11(1 downto 1) &
  n11(0 downto 0);
n14 <= unsigned(signed(n5) * signed(n12));
n15 <= n14(30 downto 30) &
  n14(29 downto 29) &
  n14(28 downto 28) &
  n14(27 downto 27) &
  n14(26 downto 26) &
  n14(25 downto 25) &
  n14(24 downto 24) &
  n14(23 downto 23) &
  n14(22 downto 22) &
  n14(21 downto 21) &
  n14(20 downto 20) &
  n14(19 downto 19) &
  n14(18 downto 18) &
  n14(17 downto 17) &
  n14(16 downto 16) &
  n14(15 downto 15);
process (clock_c) begin
  if rising_edge(clock_c) then
    if i5 = "1" then
      n16 <= "0000000000000000";
    elsif i4 = "1" then
      n16 <= n15;
    end if;
  end if;
end process;
n17 <= unsigned(signed(n6) * signed(n13));
n18 <= n17(30 downto 30) &
  n17(29 downto 29) &
  n17(28 downto 28) &
  n17(27 downto 27) &
  n17(26 downto 26) &
  n17(25 downto 25) &
  n17(24 downto 24) &
  n17(23 downto 23) &
  n17(22 downto 22) &
  n17(21 downto 21) &
  n17(20 downto 20) &
  n17(19 downto 19) &
  n17(18 downto 18) &
  n17(17 downto 17) &
  n17(16 downto 16) &
  n17(15 downto 15);
process (clock_c) begin
  if rising_edge(clock_c) then
    if i5 = "1" then
      n19 <= "0000000000000000";
    elsif i4 = "1" then
      n19 <= n18;
    end if;
  end if;
end process;
n20 <= n16 - n19;
process (clock_c) begin
  if rising_edge(clock_c) then
    if i5 = "1" then
      n21 <= "0000000000000000";
    elsif i4 = "1" then
      n21 <= n20;
    end if;
  end if;
end process;
n22 <= unsigned(signed(n5) * signed(n13));
n23 <= n22(30 downto 30) &
  n22(29 downto 29) &
  n22(28 downto 28) &
  n22(27 downto 27) &
  n22(26 downto 26) &
  n22(25 downto 25) &
  n22(24 downto 24) &
  n22(23 downto 23) &
  n22(22 downto 22) &
  n22(21 downto 21) &
  n22(20 downto 20) &
  n22(19 downto 19) &
  n22(18 downto 18) &
  n22(17 downto 17) &
  n22(16 downto 16) &
  n22(15 downto 15);
process (clock_c) begin
  if rising_edge(clock_c) then
    if i5 = "1" then
      n24 <= "0000000000000000";
    elsif i4 = "1" then
      n24 <= n23;
    end if;
  end if;
end process;
n25 <= unsigned(signed(n6) * signed(n12));
n26 <= n25(30 downto 30) &
  n25(29 downto 29) &
  n25(28 downto 28) &
  n25(27 downto 27) &
  n25(26 downto 26) &
  n25(25 downto 25) &
  n25(24 downto 24) &
  n25(23 downto 23) &
  n25(22 downto 22) &
  n25(21 downto 21) &
  n25(20 downto 20) &
  n25(19 downto 19) &
  n25(18 downto 18) &
  n25(17 downto 17) &
  n25(16 downto 16) &
  n25(15 downto 15);
process (clock_c) begin
  if rising_edge(clock_c) then
    if i5 = "1" then
      n27 <= "0000000000000000";
    elsif i4 = "1" then
      n27 <= n26;
    end if;
  end if;
end process;
n28 <= n24 + n27;
process (clock_c) begin
  if rising_edge(clock_c) then
    if i5 = "1" then
      n29 <= "0000000000000000";
    elsif i4 = "1" then
      n29 <= n28;
    end if;
  end if;
end process;
n30 <= n8 + n21;
n31 <= n10 + n29;
n32 <= n30 & n31;
process (clock_c) begin
  if rising_edge(clock_c) then
    if i5 = "1" then
      n33 <= "00000000000000000000000000000000";
    elsif i4 = "1" then
      n33 <= n32;
    end if;
  end if;
end process;
n34 <= n8 - n21;
n35 <= n10 - n29;
n36 <= n34 & n35;
process (clock_c) begin
  if rising_edge(clock_c) then
    if i5 = "1" then
      n37 <= "00000000000000000000000000000000";
    elsif i4 = "1" then
      n37 <= n36;
    end if;
  end if;
end process;
o2 <= n37;
o1 <= n33;
end architecture rtl;

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
entity cf_fft_2048_16_15 is
port (
clock_c : in std_logic;
i1 : in  unsigned(0 downto 0);
i2 : in  unsigned(31 downto 0);
i3 : in  unsigned(31 downto 0);
i4 : in  unsigned(0 downto 0);
i5 : in  unsigned(0 downto 0);
o1 : out unsigned(0 downto 0);
o2 : out unsigned(31 downto 0);
o3 : out unsigned(31 downto 0));
end entity cf_fft_2048_16_15;
architecture rtl of cf_fft_2048_16_15 is
signal n1 : unsigned(5 downto 0);
signal n2 : unsigned(63 downto 0);
signal n3 : unsigned(0 downto 0) := "0";
signal n4 : unsigned(0 downto 0) := "0";
signal n5 : unsigned(0 downto 0) := "0";
signal n6 : unsigned(0 downto 0) := "0";
signal n7 : unsigned(8 downto 0);
signal n8 : unsigned(8 downto 0) := "000000000";
signal n9 : unsigned(8 downto 0) := "000000000";
signal n10 : unsigned(8 downto 0) := "000000000";
signal n11 : unsigned(8 downto 0) := "000000000";
signal n12 : unsigned(0 downto 0);
signal n13 : unsigned(0 downto 0) := "0";
signal n14 : unsigned(0 downto 0) := "0";
signal n15 : unsigned(0 downto 0) := "0";
signal n16 : unsigned(0 downto 0) := "0";
signal n17 : unsigned(0 downto 0);
signal n18 : unsigned(1 downto 0);
signal n19 : unsigned(31 downto 0);
signal n20 : unsigned(31 downto 0);
signal n21 : unsigned(31 downto 0);
signal n22 : unsigned(31 downto 0);
signal n23 : unsigned(31 downto 0);
signal n24 : unsigned(31 downto 0);
signal s25_1 : unsigned(0 downto 0);
signal s26_1 : unsigned(31 downto 0);
signal s26_2 : unsigned(31 downto 0);
signal s27_1 : unsigned(9 downto 0);
signal s27_2 : unsigned(0 downto 0);
signal s28_1 : unsigned(0 downto 0);
signal s28_2 : unsigned(0 downto 0);
signal s28_3 : unsigned(63 downto 0);
signal s29_1 : unsigned(63 downto 0);
component cf_fft_2048_16_35 is
port (
clock_c : in std_logic;
i1 : in  unsigned(1 downto 0);
i2 : in  unsigned(0 downto 0);
i3 : in  unsigned(0 downto 0);
o1 : out unsigned(0 downto 0));
end component cf_fft_2048_16_35;
component cf_fft_2048_16_16 is
port (
clock_c : in std_logic;
i1 : in  unsigned(31 downto 0);
i2 : in  unsigned(31 downto 0);
i3 : in  unsigned(5 downto 0);
i4 : in  unsigned(0 downto 0);
i5 : in  unsigned(0 downto 0);
o1 : out unsigned(31 downto 0);
o2 : out unsigned(31 downto 0));
end component cf_fft_2048_16_16;
component cf_fft_2048_16_26 is
port (
clock_c : in std_logic;
i1 : in  unsigned(0 downto 0);
i2 : in  unsigned(0 downto 0);
i3 : in  unsigned(0 downto 0);
o1 : out unsigned(9 downto 0);
o2 : out unsigned(0 downto 0));
end component cf_fft_2048_16_26;
component cf_fft_2048_16_30 is
port (
clock_c : in std_logic;
i1 : in  unsigned(63 downto 0);
i2 : in  unsigned(0 downto 0);
i3 : in  unsigned(8 downto 0);
i4 : in  unsigned(0 downto 0);
i5 : in  unsigned(0 downto 0);
i6 : in  unsigned(0 downto 0);
o1 : out unsigned(0 downto 0);
o2 : out unsigned(0 downto 0);
o3 : out unsigned(63 downto 0));
end component cf_fft_2048_16_30;
component cf_fft_2048_16_31 is
port (
clock_c : in std_logic;
i1 : in  unsigned(63 downto 0);
i2 : in  unsigned(0 downto 0);
i3 : in  unsigned(8 downto 0);
i4 : in  unsigned(0 downto 0);
i5 : in  unsigned(0 downto 0);
i6 : in  unsigned(0 downto 0);
o1 : out unsigned(63 downto 0));
end component cf_fft_2048_16_31;
begin
n1 <= s27_1(9 downto 9) &
  s27_1(8 downto 8) &
  s27_1(7 downto 7) &
  s27_1(6 downto 6) &
  s27_1(5 downto 5) &
  s27_1(4 downto 4);
n2 <= s26_1 & s26_2;
process (clock_c) begin
  if rising_edge(clock_c) then
    if i5 = "1" then
      n3 <= "0";
    elsif i4 = "1" then
      n3 <= s27_2;
    end if;
  end if;
end process;
process (clock_c) begin
  if rising_edge(clock_c) then
    if i5 = "1" then
      n4 <= "0";
    elsif i4 = "1" then
      n4 <= n3;
    end if;
  end if;
end process;
process (clock_c) begin
  if rising_edge(clock_c) then
    if i5 = "1" then
      n5 <= "0";
    elsif i4 = "1" then
      n5 <= n4;
    end if;
  end if;
end process;
process (clock_c) begin
  if rising_edge(clock_c) then
    if i5 = "1" then
      n6 <= "0";
    elsif i4 = "1" then
      n6 <= n5;
    end if;
  end if;
end process;
n7 <= s27_1(9 downto 9) &
  s27_1(8 downto 8) &
  s27_1(7 downto 7) &
  s27_1(6 downto 6) &
  s27_1(5 downto 5) &
  s27_1(4 downto 4) &
  s27_1(3 downto 3) &
  s27_1(2 downto 2) &
  s27_1(1 downto 1);
process (clock_c) begin
  if rising_edge(clock_c) then
    if i5 = "1" then
      n8 <= "000000000";
    elsif i4 = "1" then
      n8 <= n7;
    end if;
  end if;
end process;
process (clock_c) begin
  if rising_edge(clock_c) then
    if i5 = "1" then
      n9 <= "000000000";
    elsif i4 = "1" then
      n9 <= n8;
    end if;
  end if;
end process;
process (clock_c) begin
  if rising_edge(clock_c) then
    if i5 = "1" then
      n10 <= "000000000";
    elsif i4 = "1" then
      n10 <= n9;
    end if;
  end if;
end process;
process (clock_c) begin
  if rising_edge(clock_c) then
    if i5 = "1" then
      n11 <= "000000000";
    elsif i4 = "1" then
      n11 <= n10;
    end if;
  end if;
end process;
n12 <= s27_1(0 downto 0);
process (clock_c) begin
  if rising_edge(clock_c) then
    if i5 = "1" then
      n13 <= "0";
    elsif i4 = "1" then
      n13 <= n12;
    end if;
  end if;
end process;
process (clock_c) begin
  if rising_edge(clock_c) then
    if i5 = "1" then
      n14 <= "0";
    elsif i4 = "1" then
      n14 <= n13;
    end if;
  end if;
end process;
process (clock_c) begin
  if rising_edge(clock_c) then
    if i5 = "1" then
      n15 <= "0";
    elsif i4 = "1" then
      n15 <= n14;
    end if;
  end if;
end process;
process (clock_c) begin
  if rising_edge(clock_c) then
    if i5 = "1" then
      n16 <= "0";
    elsif i4 = "1" then
      n16 <= n15;
    end if;
  end if;
end process;
n17 <= not n16;
n18 <= s28_2 & s28_1;
n19 <= s28_3(63 downto 63) &
  s28_3(62 downto 62) &
  s28_3(61 downto 61) &
  s28_3(60 downto 60) &
  s28_3(59 downto 59) &
  s28_3(58 downto 58) &
  s28_3(57 downto 57) &
  s28_3(56 downto 56) &
  s28_3(55 downto 55) &
  s28_3(54 downto 54) &
  s28_3(53 downto 53) &
  s28_3(52 downto 52) &
  s28_3(51 downto 51) &
  s28_3(50 downto 50) &
  s28_3(49 downto 49) &
  s28_3(48 downto 48) &
  s28_3(47 downto 47) &
  s28_3(46 downto 46) &
  s28_3(45 downto 45) &
  s28_3(44 downto 44) &
  s28_3(43 downto 43) &
  s28_3(42 downto 42) &
  s28_3(41 downto 41) &
  s28_3(40 downto 40) &
  s28_3(39 downto 39) &
  s28_3(38 downto 38) &
  s28_3(37 downto 37) &
  s28_3(36 downto 36) &
  s28_3(35 downto 35) &
  s28_3(34 downto 34) &
  s28_3(33 downto 33) &
  s28_3(32 downto 32);
n20 <= s28_3(31 downto 31) &
  s28_3(30 downto 30) &
  s28_3(29 downto 29) &
  s28_3(28 downto 28) &
  s28_3(27 downto 27) &
  s28_3(26 downto 26) &
  s28_3(25 downto 25) &
  s28_3(24 downto 24) &
  s28_3(23 downto 23) &
  s28_3(22 downto 22) &
  s28_3(21 downto 21) &
  s28_3(20 downto 20) &
  s28_3(19 downto 19) &
  s28_3(18 downto 18) &
  s28_3(17 downto 17) &
  s28_3(16 downto 16) &
  s28_3(15 downto 15) &
  s28_3(14 downto 14) &
  s28_3(13 downto 13) &
  s28_3(12 downto 12) &
  s28_3(11 downto 11) &
  s28_3(10 downto 10) &
  s28_3(9 downto 9) &
  s28_3(8 downto 8) &
  s28_3(7 downto 7) &
  s28_3(6 downto 6) &
  s28_3(5 downto 5) &
  s28_3(4 downto 4) &
  s28_3(3 downto 3) &
  s28_3(2 downto 2) &
  s28_3(1 downto 1) &
  s28_3(0 downto 0);
n21 <= s29_1(63 downto 63) &
  s29_1(62 downto 62) &
  s29_1(61 downto 61) &
  s29_1(60 downto 60) &
  s29_1(59 downto 59) &
  s29_1(58 downto 58) &
  s29_1(57 downto 57) &
  s29_1(56 downto 56) &
  s29_1(55 downto 55) &
  s29_1(54 downto 54) &
  s29_1(53 downto 53) &
  s29_1(52 downto 52) &
  s29_1(51 downto 51) &
  s29_1(50 downto 50) &
  s29_1(49 downto 49) &
  s29_1(48 downto 48) &
  s29_1(47 downto 47) &
  s29_1(46 downto 46) &
  s29_1(45 downto 45) &
  s29_1(44 downto 44) &
  s29_1(43 downto 43) &
  s29_1(42 downto 42) &
  s29_1(41 downto 41) &
  s29_1(40 downto 40) &
  s29_1(39 downto 39) &
  s29_1(38 downto 38) &
  s29_1(37 downto 37) &
  s29_1(36 downto 36) &
  s29_1(35 downto 35) &
  s29_1(34 downto 34) &
  s29_1(33 downto 33) &
  s29_1(32 downto 32);
n22 <= s29_1(31 downto 31) &
  s29_1(30 downto 30) &
  s29_1(29 downto 29) &
  s29_1(28 downto 28) &
  s29_1(27 downto 27) &
  s29_1(26 downto 26) &
  s29_1(25 downto 25) &
  s29_1(24 downto 24) &
  s29_1(23 downto 23) &
  s29_1(22 downto 22) &
  s29_1(21 downto 21) &
  s29_1(20 downto 20) &
  s29_1(19 downto 19) &
  s29_1(18 downto 18) &
  s29_1(17 downto 17) &
  s29_1(16 downto 16) &
  s29_1(15 downto 15) &
  s29_1(14 downto 14) &
  s29_1(13 downto 13) &
  s29_1(12 downto 12) &
  s29_1(11 downto 11) &
  s29_1(10 downto 10) &
  s29_1(9 downto 9) &
  s29_1(8 downto 8) &
  s29_1(7 downto 7) &
  s29_1(6 downto 6) &
  s29_1(5 downto 5) &
  s29_1(4 downto 4) &
  s29_1(3 downto 3) &
  s29_1(2 downto 2) &
  s29_1(1 downto 1) &
  s29_1(0 downto 0);
n23 <= n20 when s25_1 = "1" else n19;
n24 <= n22 when s25_1 = "1" else n21;
s25 : cf_fft_2048_16_35 port map (clock_c, n18, i4, i5, s25_1);
s26 : cf_fft_2048_16_16 port map (clock_c, i2, i3, n1, i4, i5, s26_1, s26_2);
s27 : cf_fft_2048_16_26 port map (clock_c, i1, i4, i5, s27_1, s27_2);
s28 : cf_fft_2048_16_30 port map (clock_c, n2, n6, n11, n17, i4, i5, s28_1, s28_2, s28_3);
s29 : cf_fft_2048_16_31 port map (clock_c, n2, n6, n11, n16, i4, i5, s29_1);
o3 <= n24;
o2 <= n23;
o1 <= s28_1;
end architecture rtl;

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
entity cf_fft_2048_16_14 is
port (
clock_c : in std_logic;
i1 : in  unsigned(31 downto 0);
i2 : in  unsigned(31 downto 0);
i3 : in  unsigned(4 downto 0);
i4 : in  unsigned(0 downto 0);
i5 : in  unsigned(0 downto 0);
o1 : out unsigned(31 downto 0);
o2 : out unsigned(31 downto 0));
end entity cf_fft_2048_16_14;
architecture rtl of cf_fft_2048_16_14 is
signal n1 : unsigned(31 downto 0) := "00000000000000000000000000000000";
signal n2 : unsigned(15 downto 0);
signal n3 : unsigned(15 downto 0);
signal n4 : unsigned(31 downto 0) := "00000000000000000000000000000000";
signal n5 : unsigned(15 downto 0);
signal n6 : unsigned(15 downto 0);
signal n7 : unsigned(15 downto 0) := "0000000000000000";
signal n8 : unsigned(15 downto 0) := "0000000000000000";
signal n9 : unsigned(15 downto 0) := "0000000000000000";
signal n10 : unsigned(15 downto 0) := "0000000000000000";
signal n11 : unsigned(31 downto 0) := "00000000000000000000000000000000";
signal n12 : unsigned(15 downto 0);
signal n13 : unsigned(15 downto 0);
signal n14 : unsigned(31 downto 0);
signal n15 : unsigned(15 downto 0);
signal n16 : unsigned(15 downto 0) := "0000000000000000";
signal n17 : unsigned(31 downto 0);
signal n18 : unsigned(15 downto 0);
signal n19 : unsigned(15 downto 0) := "0000000000000000";
signal n20 : unsigned(15 downto 0);
signal n21 : unsigned(15 downto 0) := "0000000000000000";
signal n22 : unsigned(31 downto 0);
signal n23 : unsigned(15 downto 0);
signal n24 : unsigned(15 downto 0) := "0000000000000000";
signal n25 : unsigned(31 downto 0);
signal n26 : unsigned(15 downto 0);
signal n27 : unsigned(15 downto 0) := "0000000000000000";
signal n28 : unsigned(15 downto 0);
signal n29 : unsigned(15 downto 0) := "0000000000000000";
signal n30 : unsigned(15 downto 0);
signal n31 : unsigned(15 downto 0);
signal n32 : unsigned(31 downto 0);
signal n33 : unsigned(31 downto 0) := "00000000000000000000000000000000";
signal n34 : unsigned(15 downto 0);
signal n35 : unsigned(15 downto 0);
signal n36 : unsigned(31 downto 0);
signal n37 : unsigned(31 downto 0) := "00000000000000000000000000000000";
begin
process (clock_c) begin
  if rising_edge(clock_c) then
    if i5 = "1" then
      n1 <= "00000000000000000000000000000000";
    elsif i4 = "1" then
      n1 <= i1;
    end if;
  end if;
end process;
n2 <= n1(31 downto 31) &
  n1(30 downto 30) &
  n1(29 downto 29) &
  n1(28 downto 28) &
  n1(27 downto 27) &
  n1(26 downto 26) &
  n1(25 downto 25) &
  n1(24 downto 24) &
  n1(23 downto 23) &
  n1(22 downto 22) &
  n1(21 downto 21) &
  n1(20 downto 20) &
  n1(19 downto 19) &
  n1(18 downto 18) &
  n1(17 downto 17) &
  n1(16 downto 16);
n3 <= n1(15 downto 15) &
  n1(14 downto 14) &
  n1(13 downto 13) &
  n1(12 downto 12) &
  n1(11 downto 11) &
  n1(10 downto 10) &
  n1(9 downto 9) &
  n1(8 downto 8) &
  n1(7 downto 7) &
  n1(6 downto 6) &
  n1(5 downto 5) &
  n1(4 downto 4) &
  n1(3 downto 3) &
  n1(2 downto 2) &
  n1(1 downto 1) &
  n1(0 downto 0);
process (clock_c) begin
  if rising_edge(clock_c) then
    if i5 = "1" then
      n4 <= "00000000000000000000000000000000";
    elsif i4 = "1" then
      n4 <= i2;
    end if;
  end if;
end process;
n5 <= n4(31 downto 31) &
  n4(30 downto 30) &
  n4(29 downto 29) &
  n4(28 downto 28) &
  n4(27 downto 27) &
  n4(26 downto 26) &
  n4(25 downto 25) &
  n4(24 downto 24) &
  n4(23 downto 23) &
  n4(22 downto 22) &
  n4(21 downto 21) &
  n4(20 downto 20) &
  n4(19 downto 19) &
  n4(18 downto 18) &
  n4(17 downto 17) &
  n4(16 downto 16);
n6 <= n4(15 downto 15) &
  n4(14 downto 14) &
  n4(13 downto 13) &
  n4(12 downto 12) &
  n4(11 downto 11) &
  n4(10 downto 10) &
  n4(9 downto 9) &
  n4(8 downto 8) &
  n4(7 downto 7) &
  n4(6 downto 6) &
  n4(5 downto 5) &
  n4(4 downto 4) &
  n4(3 downto 3) &
  n4(2 downto 2) &
  n4(1 downto 1) &
  n4(0 downto 0);
process (clock_c) begin
  if rising_edge(clock_c) then
    if i5 = "1" then
      n7 <= "0000000000000000";
    elsif i4 = "1" then
      n7 <= n2;
    end if;
  end if;
end process;
process (clock_c) begin
  if rising_edge(clock_c) then
    if i5 = "1" then
      n8 <= "0000000000000000";
    elsif i4 = "1" then
      n8 <= n7;
    end if;
  end if;
end process;
process (clock_c) begin
  if rising_edge(clock_c) then
    if i5 = "1" then
      n9 <= "0000000000000000";
    elsif i4 = "1" then
      n9 <= n3;
    end if;
  end if;
end process;
process (clock_c) begin
  if rising_edge(clock_c) then
    if i5 = "1" then
      n10 <= "0000000000000000";
    elsif i4 = "1" then
      n10 <= n9;
    end if;
  end if;
end process;
process (clock_c) begin
  if rising_edge(clock_c) then 
    if i4 = "1" then
      case i3 is
        when "00000" => n11 <= "01111111111111110000000000000000";
        when "00001" => n11 <= "01111111011000101111001101110100";
        when "00010" => n11 <= "01111101100010101110011100000111";
        when "00011" => n11 <= "01111010011111011101101011010111";
        when "00100" => n11 <= "01110110010000011100111100000100";
        when "00101" => n11 <= "01110000111000101100001110101001";
        when "00110" => n11 <= "01101010011011011011100011100011";
        when "00111" => n11 <= "01100010111100101010111011001100";
        when "01000" => n11 <= "01011010100000101010010101111101";
        when "01001" => n11 <= "01010001001100111001110100001101";
        when "01010" => n11 <= "01000111000111001001010110010010";
        when "01011" => n11 <= "00111100010101101000111100011101";
        when "01100" => n11 <= "00110000111110111000100110111110";
        when "01101" => n11 <= "00100101001010001000010110000010";
        when "01110" => n11 <= "00011000111110001000001001110101";
        when "01111" => n11 <= "00001100100010111000000010011101";
        when "10000" => n11 <= "00000000000000001000000000000000";
        when "10001" => n11 <= "11110011011101001000000010011101";
        when "10010" => n11 <= "11100111000001111000001001110101";
        when "10011" => n11 <= "11011010110101111000010110000010";
        when "10100" => n11 <= "11001111000001001000100110111110";
        when "10101" => n11 <= "11000011101010011000111100011101";
        when "10110" => n11 <= "10111000111000111001010110010010";
        when "10111" => n11 <= "10101110110011001001110100001101";
        when "11000" => n11 <= "10100101011111011010010101111101";
        when "11001" => n11 <= "10011101000011011010111011001100";
        when "11010" => n11 <= "10010101100100101011100011100011";
        when "11011" => n11 <= "10001111000111011100001110101001";
        when "11100" => n11 <= "10001001101111101100111100000100";
        when "11101" => n11 <= "10000101100000101101101011010111";
        when "11110" => n11 <= "10000010011101011110011100000111";
        when "11111" => n11 <= "10000000100111011111001101110100";
        when others => n11 <= "XXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX";
      end case;
    end if;
  end if;
end process;
n12 <= n11(31 downto 31) &
  n11(30 downto 30) &
  n11(29 downto 29) &
  n11(28 downto 28) &
  n11(27 downto 27) &
  n11(26 downto 26) &
  n11(25 downto 25) &
  n11(24 downto 24) &
  n11(23 downto 23) &
  n11(22 downto 22) &
  n11(21 downto 21) &
  n11(20 downto 20) &
  n11(19 downto 19) &
  n11(18 downto 18) &
  n11(17 downto 17) &
  n11(16 downto 16);
n13 <= n11(15 downto 15) &
  n11(14 downto 14) &
  n11(13 downto 13) &
  n11(12 downto 12) &
  n11(11 downto 11) &
  n11(10 downto 10) &
  n11(9 downto 9) &
  n11(8 downto 8) &
  n11(7 downto 7) &
  n11(6 downto 6) &
  n11(5 downto 5) &
  n11(4 downto 4) &
  n11(3 downto 3) &
  n11(2 downto 2) &
  n11(1 downto 1) &
  n11(0 downto 0);
n14 <= unsigned(signed(n5) * signed(n12));
n15 <= n14(30 downto 30) &
  n14(29 downto 29) &
  n14(28 downto 28) &
  n14(27 downto 27) &
  n14(26 downto 26) &
  n14(25 downto 25) &
  n14(24 downto 24) &
  n14(23 downto 23) &
  n14(22 downto 22) &
  n14(21 downto 21) &
  n14(20 downto 20) &
  n14(19 downto 19) &
  n14(18 downto 18) &
  n14(17 downto 17) &
  n14(16 downto 16) &
  n14(15 downto 15);
process (clock_c) begin
  if rising_edge(clock_c) then
    if i5 = "1" then
      n16 <= "0000000000000000";
    elsif i4 = "1" then
      n16 <= n15;
    end if;
  end if;
end process;
n17 <= unsigned(signed(n6) * signed(n13));
n18 <= n17(30 downto 30) &
  n17(29 downto 29) &
  n17(28 downto 28) &
  n17(27 downto 27) &
  n17(26 downto 26) &
  n17(25 downto 25) &
  n17(24 downto 24) &
  n17(23 downto 23) &
  n17(22 downto 22) &
  n17(21 downto 21) &
  n17(20 downto 20) &
  n17(19 downto 19) &
  n17(18 downto 18) &
  n17(17 downto 17) &
  n17(16 downto 16) &
  n17(15 downto 15);
process (clock_c) begin
  if rising_edge(clock_c) then
    if i5 = "1" then
      n19 <= "0000000000000000";
    elsif i4 = "1" then
      n19 <= n18;
    end if;
  end if;
end process;
n20 <= n16 - n19;
process (clock_c) begin
  if rising_edge(clock_c) then
    if i5 = "1" then
      n21 <= "0000000000000000";
    elsif i4 = "1" then
      n21 <= n20;
    end if;
  end if;
end process;
n22 <= unsigned(signed(n5) * signed(n13));
n23 <= n22(30 downto 30) &
  n22(29 downto 29) &
  n22(28 downto 28) &
  n22(27 downto 27) &
  n22(26 downto 26) &
  n22(25 downto 25) &
  n22(24 downto 24) &
  n22(23 downto 23) &
  n22(22 downto 22) &
  n22(21 downto 21) &
  n22(20 downto 20) &
  n22(19 downto 19) &
  n22(18 downto 18) &
  n22(17 downto 17) &
  n22(16 downto 16) &
  n22(15 downto 15);
process (clock_c) begin
  if rising_edge(clock_c) then
    if i5 = "1" then
      n24 <= "0000000000000000";
    elsif i4 = "1" then
      n24 <= n23;
    end if;
  end if;
end process;
n25 <= unsigned(signed(n6) * signed(n12));
n26 <= n25(30 downto 30) &
  n25(29 downto 29) &
  n25(28 downto 28) &
  n25(27 downto 27) &
  n25(26 downto 26) &
  n25(25 downto 25) &
  n25(24 downto 24) &
  n25(23 downto 23) &
  n25(22 downto 22) &
  n25(21 downto 21) &
  n25(20 downto 20) &
  n25(19 downto 19) &
  n25(18 downto 18) &
  n25(17 downto 17) &
  n25(16 downto 16) &
  n25(15 downto 15);
process (clock_c) begin
  if rising_edge(clock_c) then
    if i5 = "1" then
      n27 <= "0000000000000000";
    elsif i4 = "1" then
      n27 <= n26;
    end if;
  end if;
end process;
n28 <= n24 + n27;
process (clock_c) begin
  if rising_edge(clock_c) then
    if i5 = "1" then
      n29 <= "0000000000000000";
    elsif i4 = "1" then
      n29 <= n28;
    end if;
  end if;
end process;
n30 <= n8 + n21;
n31 <= n10 + n29;
n32 <= n30 & n31;
process (clock_c) begin
  if rising_edge(clock_c) then
    if i5 = "1" then
      n33 <= "00000000000000000000000000000000";
    elsif i4 = "1" then
      n33 <= n32;
    end if;
  end if;
end process;
n34 <= n8 - n21;
n35 <= n10 - n29;
n36 <= n34 & n35;
process (clock_c) begin
  if rising_edge(clock_c) then
    if i5 = "1" then
      n37 <= "00000000000000000000000000000000";
    elsif i4 = "1" then
      n37 <= n36;
    end if;
  end if;
end process;
o2 <= n37;
o1 <= n33;
end architecture rtl;

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
entity cf_fft_2048_16_13 is
port (
clock_c : in std_logic;
i1 : in  unsigned(0 downto 0);
i2 : in  unsigned(31 downto 0);
i3 : in  unsigned(31 downto 0);
i4 : in  unsigned(0 downto 0);
i5 : in  unsigned(0 downto 0);
o1 : out unsigned(0 downto 0);
o2 : out unsigned(31 downto 0);
o3 : out unsigned(31 downto 0));
end entity cf_fft_2048_16_13;
architecture rtl of cf_fft_2048_16_13 is
signal n1 : unsigned(4 downto 0);
signal n2 : unsigned(63 downto 0);
signal n3 : unsigned(0 downto 0) := "0";
signal n4 : unsigned(0 downto 0) := "0";
signal n5 : unsigned(0 downto 0) := "0";
signal n6 : unsigned(0 downto 0) := "0";
signal n7 : unsigned(8 downto 0);
signal n8 : unsigned(8 downto 0) := "000000000";
signal n9 : unsigned(8 downto 0) := "000000000";
signal n10 : unsigned(8 downto 0) := "000000000";
signal n11 : unsigned(8 downto 0) := "000000000";
signal n12 : unsigned(0 downto 0);
signal n13 : unsigned(0 downto 0) := "0";
signal n14 : unsigned(0 downto 0) := "0";
signal n15 : unsigned(0 downto 0) := "0";
signal n16 : unsigned(0 downto 0) := "0";
signal n17 : unsigned(0 downto 0);
signal n18 : unsigned(1 downto 0);
signal n19 : unsigned(31 downto 0);
signal n20 : unsigned(31 downto 0);
signal n21 : unsigned(31 downto 0);
signal n22 : unsigned(31 downto 0);
signal n23 : unsigned(31 downto 0);
signal n24 : unsigned(31 downto 0);
signal s25_1 : unsigned(0 downto 0);
signal s26_1 : unsigned(31 downto 0);
signal s26_2 : unsigned(31 downto 0);
signal s27_1 : unsigned(9 downto 0);
signal s27_2 : unsigned(0 downto 0);
signal s28_1 : unsigned(0 downto 0);
signal s28_2 : unsigned(0 downto 0);
signal s28_3 : unsigned(63 downto 0);
signal s29_1 : unsigned(63 downto 0);
component cf_fft_2048_16_35 is
port (
clock_c : in std_logic;
i1 : in  unsigned(1 downto 0);
i2 : in  unsigned(0 downto 0);
i3 : in  unsigned(0 downto 0);
o1 : out unsigned(0 downto 0));
end component cf_fft_2048_16_35;
component cf_fft_2048_16_14 is
port (
clock_c : in std_logic;
i1 : in  unsigned(31 downto 0);
i2 : in  unsigned(31 downto 0);
i3 : in  unsigned(4 downto 0);
i4 : in  unsigned(0 downto 0);
i5 : in  unsigned(0 downto 0);
o1 : out unsigned(31 downto 0);
o2 : out unsigned(31 downto 0));
end component cf_fft_2048_16_14;
component cf_fft_2048_16_26 is
port (
clock_c : in std_logic;
i1 : in  unsigned(0 downto 0);
i2 : in  unsigned(0 downto 0);
i3 : in  unsigned(0 downto 0);
o1 : out unsigned(9 downto 0);
o2 : out unsigned(0 downto 0));
end component cf_fft_2048_16_26;
component cf_fft_2048_16_30 is
port (
clock_c : in std_logic;
i1 : in  unsigned(63 downto 0);
i2 : in  unsigned(0 downto 0);
i3 : in  unsigned(8 downto 0);
i4 : in  unsigned(0 downto 0);
i5 : in  unsigned(0 downto 0);
i6 : in  unsigned(0 downto 0);
o1 : out unsigned(0 downto 0);
o2 : out unsigned(0 downto 0);
o3 : out unsigned(63 downto 0));
end component cf_fft_2048_16_30;
component cf_fft_2048_16_31 is
port (
clock_c : in std_logic;
i1 : in  unsigned(63 downto 0);
i2 : in  unsigned(0 downto 0);
i3 : in  unsigned(8 downto 0);
i4 : in  unsigned(0 downto 0);
i5 : in  unsigned(0 downto 0);
i6 : in  unsigned(0 downto 0);
o1 : out unsigned(63 downto 0));
end component cf_fft_2048_16_31;
begin
n1 <= s27_1(9 downto 9) &
  s27_1(8 downto 8) &
  s27_1(7 downto 7) &
  s27_1(6 downto 6) &
  s27_1(5 downto 5);
n2 <= s26_1 & s26_2;
process (clock_c) begin
  if rising_edge(clock_c) then
    if i5 = "1" then
      n3 <= "0";
    elsif i4 = "1" then
      n3 <= s27_2;
    end if;
  end if;
end process;
process (clock_c) begin
  if rising_edge(clock_c) then
    if i5 = "1" then
      n4 <= "0";
    elsif i4 = "1" then
      n4 <= n3;
    end if;
  end if;
end process;
process (clock_c) begin
  if rising_edge(clock_c) then
    if i5 = "1" then
      n5 <= "0";
    elsif i4 = "1" then
      n5 <= n4;
    end if;
  end if;
end process;
process (clock_c) begin
  if rising_edge(clock_c) then
    if i5 = "1" then
      n6 <= "0";
    elsif i4 = "1" then
      n6 <= n5;
    end if;
  end if;
end process;
n7 <= s27_1(9 downto 9) &
  s27_1(8 downto 8) &
  s27_1(7 downto 7) &
  s27_1(6 downto 6) &
  s27_1(5 downto 5) &
  s27_1(4 downto 4) &
  s27_1(3 downto 3) &
  s27_1(2 downto 2) &
  s27_1(1 downto 1);
process (clock_c) begin
  if rising_edge(clock_c) then
    if i5 = "1" then
      n8 <= "000000000";
    elsif i4 = "1" then
      n8 <= n7;
    end if;
  end if;
end process;
process (clock_c) begin
  if rising_edge(clock_c) then
    if i5 = "1" then
      n9 <= "000000000";
    elsif i4 = "1" then
      n9 <= n8;
    end if;
  end if;
end process;
process (clock_c) begin
  if rising_edge(clock_c) then
    if i5 = "1" then
      n10 <= "000000000";
    elsif i4 = "1" then
      n10 <= n9;
    end if;
  end if;
end process;
process (clock_c) begin
  if rising_edge(clock_c) then
    if i5 = "1" then
      n11 <= "000000000";
    elsif i4 = "1" then
      n11 <= n10;
    end if;
  end if;
end process;
n12 <= s27_1(0 downto 0);
process (clock_c) begin
  if rising_edge(clock_c) then
    if i5 = "1" then
      n13 <= "0";
    elsif i4 = "1" then
      n13 <= n12;
    end if;
  end if;
end process;
process (clock_c) begin
  if rising_edge(clock_c) then
    if i5 = "1" then
      n14 <= "0";
    elsif i4 = "1" then
      n14 <= n13;
    end if;
  end if;
end process;
process (clock_c) begin
  if rising_edge(clock_c) then
    if i5 = "1" then
      n15 <= "0";
    elsif i4 = "1" then
      n15 <= n14;
    end if;
  end if;
end process;
process (clock_c) begin
  if rising_edge(clock_c) then
    if i5 = "1" then
      n16 <= "0";
    elsif i4 = "1" then
      n16 <= n15;
    end if;
  end if;
end process;
n17 <= not n16;
n18 <= s28_2 & s28_1;
n19 <= s28_3(63 downto 63) &
  s28_3(62 downto 62) &
  s28_3(61 downto 61) &
  s28_3(60 downto 60) &
  s28_3(59 downto 59) &
  s28_3(58 downto 58) &
  s28_3(57 downto 57) &
  s28_3(56 downto 56) &
  s28_3(55 downto 55) &
  s28_3(54 downto 54) &
  s28_3(53 downto 53) &
  s28_3(52 downto 52) &
  s28_3(51 downto 51) &
  s28_3(50 downto 50) &
  s28_3(49 downto 49) &
  s28_3(48 downto 48) &
  s28_3(47 downto 47) &
  s28_3(46 downto 46) &
  s28_3(45 downto 45) &
  s28_3(44 downto 44) &
  s28_3(43 downto 43) &
  s28_3(42 downto 42) &
  s28_3(41 downto 41) &
  s28_3(40 downto 40) &
  s28_3(39 downto 39) &
  s28_3(38 downto 38) &
  s28_3(37 downto 37) &
  s28_3(36 downto 36) &
  s28_3(35 downto 35) &
  s28_3(34 downto 34) &
  s28_3(33 downto 33) &
  s28_3(32 downto 32);
n20 <= s28_3(31 downto 31) &
  s28_3(30 downto 30) &
  s28_3(29 downto 29) &
  s28_3(28 downto 28) &
  s28_3(27 downto 27) &
  s28_3(26 downto 26) &
  s28_3(25 downto 25) &
  s28_3(24 downto 24) &
  s28_3(23 downto 23) &
  s28_3(22 downto 22) &
  s28_3(21 downto 21) &
  s28_3(20 downto 20) &
  s28_3(19 downto 19) &
  s28_3(18 downto 18) &
  s28_3(17 downto 17) &
  s28_3(16 downto 16) &
  s28_3(15 downto 15) &
  s28_3(14 downto 14) &
  s28_3(13 downto 13) &
  s28_3(12 downto 12) &
  s28_3(11 downto 11) &
  s28_3(10 downto 10) &
  s28_3(9 downto 9) &
  s28_3(8 downto 8) &
  s28_3(7 downto 7) &
  s28_3(6 downto 6) &
  s28_3(5 downto 5) &
  s28_3(4 downto 4) &
  s28_3(3 downto 3) &
  s28_3(2 downto 2) &
  s28_3(1 downto 1) &
  s28_3(0 downto 0);
n21 <= s29_1(63 downto 63) &
  s29_1(62 downto 62) &
  s29_1(61 downto 61) &
  s29_1(60 downto 60) &
  s29_1(59 downto 59) &
  s29_1(58 downto 58) &
  s29_1(57 downto 57) &
  s29_1(56 downto 56) &
  s29_1(55 downto 55) &
  s29_1(54 downto 54) &
  s29_1(53 downto 53) &
  s29_1(52 downto 52) &
  s29_1(51 downto 51) &
  s29_1(50 downto 50) &
  s29_1(49 downto 49) &
  s29_1(48 downto 48) &
  s29_1(47 downto 47) &
  s29_1(46 downto 46) &
  s29_1(45 downto 45) &
  s29_1(44 downto 44) &
  s29_1(43 downto 43) &
  s29_1(42 downto 42) &
  s29_1(41 downto 41) &
  s29_1(40 downto 40) &
  s29_1(39 downto 39) &
  s29_1(38 downto 38) &
  s29_1(37 downto 37) &
  s29_1(36 downto 36) &
  s29_1(35 downto 35) &
  s29_1(34 downto 34) &
  s29_1(33 downto 33) &
  s29_1(32 downto 32);
n22 <= s29_1(31 downto 31) &
  s29_1(30 downto 30) &
  s29_1(29 downto 29) &
  s29_1(28 downto 28) &
  s29_1(27 downto 27) &
  s29_1(26 downto 26) &
  s29_1(25 downto 25) &
  s29_1(24 downto 24) &
  s29_1(23 downto 23) &
  s29_1(22 downto 22) &
  s29_1(21 downto 21) &
  s29_1(20 downto 20) &
  s29_1(19 downto 19) &
  s29_1(18 downto 18) &
  s29_1(17 downto 17) &
  s29_1(16 downto 16) &
  s29_1(15 downto 15) &
  s29_1(14 downto 14) &
  s29_1(13 downto 13) &
  s29_1(12 downto 12) &
  s29_1(11 downto 11) &
  s29_1(10 downto 10) &
  s29_1(9 downto 9) &
  s29_1(8 downto 8) &
  s29_1(7 downto 7) &
  s29_1(6 downto 6) &
  s29_1(5 downto 5) &
  s29_1(4 downto 4) &
  s29_1(3 downto 3) &
  s29_1(2 downto 2) &
  s29_1(1 downto 1) &
  s29_1(0 downto 0);
n23 <= n20 when s25_1 = "1" else n19;
n24 <= n22 when s25_1 = "1" else n21;
s25 : cf_fft_2048_16_35 port map (clock_c, n18, i4, i5, s25_1);
s26 : cf_fft_2048_16_14 port map (clock_c, i2, i3, n1, i4, i5, s26_1, s26_2);
s27 : cf_fft_2048_16_26 port map (clock_c, i1, i4, i5, s27_1, s27_2);
s28 : cf_fft_2048_16_30 port map (clock_c, n2, n6, n11, n17, i4, i5, s28_1, s28_2, s28_3);
s29 : cf_fft_2048_16_31 port map (clock_c, n2, n6, n11, n16, i4, i5, s29_1);
o3 <= n24;
o2 <= n23;
o1 <= s28_1;
end architecture rtl;

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
entity cf_fft_2048_16_12 is
port (
clock_c : in std_logic;
i1 : in  unsigned(31 downto 0);
i2 : in  unsigned(31 downto 0);
i3 : in  unsigned(3 downto 0);
i4 : in  unsigned(0 downto 0);
i5 : in  unsigned(0 downto 0);
o1 : out unsigned(31 downto 0);
o2 : out unsigned(31 downto 0));
end entity cf_fft_2048_16_12;
architecture rtl of cf_fft_2048_16_12 is
signal n1 : unsigned(31 downto 0) := "00000000000000000000000000000000";
signal n2 : unsigned(15 downto 0);
signal n3 : unsigned(15 downto 0);
signal n4 : unsigned(31 downto 0) := "00000000000000000000000000000000";
signal n5 : unsigned(15 downto 0);
signal n6 : unsigned(15 downto 0);
signal n7 : unsigned(15 downto 0) := "0000000000000000";
signal n8 : unsigned(15 downto 0) := "0000000000000000";
signal n9 : unsigned(15 downto 0) := "0000000000000000";
signal n10 : unsigned(15 downto 0) := "0000000000000000";
signal n11 : unsigned(31 downto 0) := "00000000000000000000000000000000";
signal n12 : unsigned(15 downto 0);
signal n13 : unsigned(15 downto 0);
signal n14 : unsigned(31 downto 0);
signal n15 : unsigned(15 downto 0);
signal n16 : unsigned(15 downto 0) := "0000000000000000";
signal n17 : unsigned(31 downto 0);
signal n18 : unsigned(15 downto 0);
signal n19 : unsigned(15 downto 0) := "0000000000000000";
signal n20 : unsigned(15 downto 0);
signal n21 : unsigned(15 downto 0) := "0000000000000000";
signal n22 : unsigned(31 downto 0);
signal n23 : unsigned(15 downto 0);
signal n24 : unsigned(15 downto 0) := "0000000000000000";
signal n25 : unsigned(31 downto 0);
signal n26 : unsigned(15 downto 0);
signal n27 : unsigned(15 downto 0) := "0000000000000000";
signal n28 : unsigned(15 downto 0);
signal n29 : unsigned(15 downto 0) := "0000000000000000";
signal n30 : unsigned(15 downto 0);
signal n31 : unsigned(15 downto 0);
signal n32 : unsigned(31 downto 0);
signal n33 : unsigned(31 downto 0) := "00000000000000000000000000000000";
signal n34 : unsigned(15 downto 0);
signal n35 : unsigned(15 downto 0);
signal n36 : unsigned(31 downto 0);
signal n37 : unsigned(31 downto 0) := "00000000000000000000000000000000";
begin
process (clock_c) begin
  if rising_edge(clock_c) then
    if i5 = "1" then
      n1 <= "00000000000000000000000000000000";
    elsif i4 = "1" then
      n1 <= i1;
    end if;
  end if;
end process;
n2 <= n1(31 downto 31) &
  n1(30 downto 30) &
  n1(29 downto 29) &
  n1(28 downto 28) &
  n1(27 downto 27) &
  n1(26 downto 26) &
  n1(25 downto 25) &
  n1(24 downto 24) &
  n1(23 downto 23) &
  n1(22 downto 22) &
  n1(21 downto 21) &
  n1(20 downto 20) &
  n1(19 downto 19) &
  n1(18 downto 18) &
  n1(17 downto 17) &
  n1(16 downto 16);
n3 <= n1(15 downto 15) &
  n1(14 downto 14) &
  n1(13 downto 13) &
  n1(12 downto 12) &
  n1(11 downto 11) &
  n1(10 downto 10) &
  n1(9 downto 9) &
  n1(8 downto 8) &
  n1(7 downto 7) &
  n1(6 downto 6) &
  n1(5 downto 5) &
  n1(4 downto 4) &
  n1(3 downto 3) &
  n1(2 downto 2) &
  n1(1 downto 1) &
  n1(0 downto 0);
process (clock_c) begin
  if rising_edge(clock_c) then
    if i5 = "1" then
      n4 <= "00000000000000000000000000000000";
    elsif i4 = "1" then
      n4 <= i2;
    end if;
  end if;
end process;
n5 <= n4(31 downto 31) &
  n4(30 downto 30) &
  n4(29 downto 29) &
  n4(28 downto 28) &
  n4(27 downto 27) &
  n4(26 downto 26) &
  n4(25 downto 25) &
  n4(24 downto 24) &
  n4(23 downto 23) &
  n4(22 downto 22) &
  n4(21 downto 21) &
  n4(20 downto 20) &
  n4(19 downto 19) &
  n4(18 downto 18) &
  n4(17 downto 17) &
  n4(16 downto 16);
n6 <= n4(15 downto 15) &
  n4(14 downto 14) &
  n4(13 downto 13) &
  n4(12 downto 12) &
  n4(11 downto 11) &
  n4(10 downto 10) &
  n4(9 downto 9) &
  n4(8 downto 8) &
  n4(7 downto 7) &
  n4(6 downto 6) &
  n4(5 downto 5) &
  n4(4 downto 4) &
  n4(3 downto 3) &
  n4(2 downto 2) &
  n4(1 downto 1) &
  n4(0 downto 0);
process (clock_c) begin
  if rising_edge(clock_c) then
    if i5 = "1" then
      n7 <= "0000000000000000";
    elsif i4 = "1" then
      n7 <= n2;
    end if;
  end if;
end process;
process (clock_c) begin
  if rising_edge(clock_c) then
    if i5 = "1" then
      n8 <= "0000000000000000";
    elsif i4 = "1" then
      n8 <= n7;
    end if;
  end if;
end process;
process (clock_c) begin
  if rising_edge(clock_c) then
    if i5 = "1" then
      n9 <= "0000000000000000";
    elsif i4 = "1" then
      n9 <= n3;
    end if;
  end if;
end process;
process (clock_c) begin
  if rising_edge(clock_c) then
    if i5 = "1" then
      n10 <= "0000000000000000";
    elsif i4 = "1" then
      n10 <= n9;
    end if;
  end if;
end process;
process (clock_c) begin
  if rising_edge(clock_c) then 
    if i4 = "1" then
      case i3 is
        when "0000" => n11 <= "01111111111111110000000000000000";
        when "0001" => n11 <= "01111101100010101110011100000111";
        when "0010" => n11 <= "01110110010000011100111100000100";
        when "0011" => n11 <= "01101010011011011011100011100011";
        when "0100" => n11 <= "01011010100000101010010101111101";
        when "0101" => n11 <= "01000111000111001001010110010010";
        when "0110" => n11 <= "00110000111110111000100110111110";
        when "0111" => n11 <= "00011000111110001000001001110101";
        when "1000" => n11 <= "00000000000000001000000000000000";
        when "1001" => n11 <= "11100111000001111000001001110101";
        when "1010" => n11 <= "11001111000001001000100110111110";
        when "1011" => n11 <= "10111000111000111001010110010010";
        when "1100" => n11 <= "10100101011111011010010101111101";
        when "1101" => n11 <= "10010101100100101011100011100011";
        when "1110" => n11 <= "10001001101111101100111100000100";
        when "1111" => n11 <= "10000010011101011110011100000111";
        when others => n11 <= "XXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX";
      end case;
    end if;
  end if;
end process;
n12 <= n11(31 downto 31) &
  n11(30 downto 30) &
  n11(29 downto 29) &
  n11(28 downto 28) &
  n11(27 downto 27) &
  n11(26 downto 26) &
  n11(25 downto 25) &
  n11(24 downto 24) &
  n11(23 downto 23) &
  n11(22 downto 22) &
  n11(21 downto 21) &
  n11(20 downto 20) &
  n11(19 downto 19) &
  n11(18 downto 18) &
  n11(17 downto 17) &
  n11(16 downto 16);
n13 <= n11(15 downto 15) &
  n11(14 downto 14) &
  n11(13 downto 13) &
  n11(12 downto 12) &
  n11(11 downto 11) &
  n11(10 downto 10) &
  n11(9 downto 9) &
  n11(8 downto 8) &
  n11(7 downto 7) &
  n11(6 downto 6) &
  n11(5 downto 5) &
  n11(4 downto 4) &
  n11(3 downto 3) &
  n11(2 downto 2) &
  n11(1 downto 1) &
  n11(0 downto 0);
n14 <= unsigned(signed(n5) * signed(n12));
n15 <= n14(30 downto 30) &
  n14(29 downto 29) &
  n14(28 downto 28) &
  n14(27 downto 27) &
  n14(26 downto 26) &
  n14(25 downto 25) &
  n14(24 downto 24) &
  n14(23 downto 23) &
  n14(22 downto 22) &
  n14(21 downto 21) &
  n14(20 downto 20) &
  n14(19 downto 19) &
  n14(18 downto 18) &
  n14(17 downto 17) &
  n14(16 downto 16) &
  n14(15 downto 15);
process (clock_c) begin
  if rising_edge(clock_c) then
    if i5 = "1" then
      n16 <= "0000000000000000";
    elsif i4 = "1" then
      n16 <= n15;
    end if;
  end if;
end process;
n17 <= unsigned(signed(n6) * signed(n13));
n18 <= n17(30 downto 30) &
  n17(29 downto 29) &
  n17(28 downto 28) &
  n17(27 downto 27) &
  n17(26 downto 26) &
  n17(25 downto 25) &
  n17(24 downto 24) &
  n17(23 downto 23) &
  n17(22 downto 22) &
  n17(21 downto 21) &
  n17(20 downto 20) &
  n17(19 downto 19) &
  n17(18 downto 18) &
  n17(17 downto 17) &
  n17(16 downto 16) &
  n17(15 downto 15);
process (clock_c) begin
  if rising_edge(clock_c) then
    if i5 = "1" then
      n19 <= "0000000000000000";
    elsif i4 = "1" then
      n19 <= n18;
    end if;
  end if;
end process;
n20 <= n16 - n19;
process (clock_c) begin
  if rising_edge(clock_c) then
    if i5 = "1" then
      n21 <= "0000000000000000";
    elsif i4 = "1" then
      n21 <= n20;
    end if;
  end if;
end process;
n22 <= unsigned(signed(n5) * signed(n13));
n23 <= n22(30 downto 30) &
  n22(29 downto 29) &
  n22(28 downto 28) &
  n22(27 downto 27) &
  n22(26 downto 26) &
  n22(25 downto 25) &
  n22(24 downto 24) &
  n22(23 downto 23) &
  n22(22 downto 22) &
  n22(21 downto 21) &
  n22(20 downto 20) &
  n22(19 downto 19) &
  n22(18 downto 18) &
  n22(17 downto 17) &
  n22(16 downto 16) &
  n22(15 downto 15);
process (clock_c) begin
  if rising_edge(clock_c) then
    if i5 = "1" then
      n24 <= "0000000000000000";
    elsif i4 = "1" then
      n24 <= n23;
    end if;
  end if;
end process;
n25 <= unsigned(signed(n6) * signed(n12));
n26 <= n25(30 downto 30) &
  n25(29 downto 29) &
  n25(28 downto 28) &
  n25(27 downto 27) &
  n25(26 downto 26) &
  n25(25 downto 25) &
  n25(24 downto 24) &
  n25(23 downto 23) &
  n25(22 downto 22) &
  n25(21 downto 21) &
  n25(20 downto 20) &
  n25(19 downto 19) &
  n25(18 downto 18) &
  n25(17 downto 17) &
  n25(16 downto 16) &
  n25(15 downto 15);
process (clock_c) begin
  if rising_edge(clock_c) then
    if i5 = "1" then
      n27 <= "0000000000000000";
    elsif i4 = "1" then
      n27 <= n26;
    end if;
  end if;
end process;
n28 <= n24 + n27;
process (clock_c) begin
  if rising_edge(clock_c) then
    if i5 = "1" then
      n29 <= "0000000000000000";
    elsif i4 = "1" then
      n29 <= n28;
    end if;
  end if;
end process;
n30 <= n8 + n21;
n31 <= n10 + n29;
n32 <= n30 & n31;
process (clock_c) begin
  if rising_edge(clock_c) then
    if i5 = "1" then
      n33 <= "00000000000000000000000000000000";
    elsif i4 = "1" then
      n33 <= n32;
    end if;
  end if;
end process;
n34 <= n8 - n21;
n35 <= n10 - n29;
n36 <= n34 & n35;
process (clock_c) begin
  if rising_edge(clock_c) then
    if i5 = "1" then
      n37 <= "00000000000000000000000000000000";
    elsif i4 = "1" then
      n37 <= n36;
    end if;
  end if;
end process;
o2 <= n37;
o1 <= n33;
end architecture rtl;

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
entity cf_fft_2048_16_11 is
port (
clock_c : in std_logic;
i1 : in  unsigned(0 downto 0);
i2 : in  unsigned(31 downto 0);
i3 : in  unsigned(31 downto 0);
i4 : in  unsigned(0 downto 0);
i5 : in  unsigned(0 downto 0);
o1 : out unsigned(0 downto 0);
o2 : out unsigned(31 downto 0);
o3 : out unsigned(31 downto 0));
end entity cf_fft_2048_16_11;
architecture rtl of cf_fft_2048_16_11 is
signal n1 : unsigned(3 downto 0);
signal n2 : unsigned(63 downto 0);
signal n3 : unsigned(0 downto 0) := "0";
signal n4 : unsigned(0 downto 0) := "0";
signal n5 : unsigned(0 downto 0) := "0";
signal n6 : unsigned(0 downto 0) := "0";
signal n7 : unsigned(8 downto 0);
signal n8 : unsigned(8 downto 0) := "000000000";
signal n9 : unsigned(8 downto 0) := "000000000";
signal n10 : unsigned(8 downto 0) := "000000000";
signal n11 : unsigned(8 downto 0) := "000000000";
signal n12 : unsigned(0 downto 0);
signal n13 : unsigned(0 downto 0) := "0";
signal n14 : unsigned(0 downto 0) := "0";
signal n15 : unsigned(0 downto 0) := "0";
signal n16 : unsigned(0 downto 0) := "0";
signal n17 : unsigned(0 downto 0);
signal n18 : unsigned(1 downto 0);
signal n19 : unsigned(31 downto 0);
signal n20 : unsigned(31 downto 0);
signal n21 : unsigned(31 downto 0);
signal n22 : unsigned(31 downto 0);
signal n23 : unsigned(31 downto 0);
signal n24 : unsigned(31 downto 0);
signal s25_1 : unsigned(0 downto 0);
signal s26_1 : unsigned(31 downto 0);
signal s26_2 : unsigned(31 downto 0);
signal s27_1 : unsigned(9 downto 0);
signal s27_2 : unsigned(0 downto 0);
signal s28_1 : unsigned(0 downto 0);
signal s28_2 : unsigned(0 downto 0);
signal s28_3 : unsigned(63 downto 0);
signal s29_1 : unsigned(63 downto 0);
component cf_fft_2048_16_35 is
port (
clock_c : in std_logic;
i1 : in  unsigned(1 downto 0);
i2 : in  unsigned(0 downto 0);
i3 : in  unsigned(0 downto 0);
o1 : out unsigned(0 downto 0));
end component cf_fft_2048_16_35;
component cf_fft_2048_16_12 is
port (
clock_c : in std_logic;
i1 : in  unsigned(31 downto 0);
i2 : in  unsigned(31 downto 0);
i3 : in  unsigned(3 downto 0);
i4 : in  unsigned(0 downto 0);
i5 : in  unsigned(0 downto 0);
o1 : out unsigned(31 downto 0);
o2 : out unsigned(31 downto 0));
end component cf_fft_2048_16_12;
component cf_fft_2048_16_26 is
port (
clock_c : in std_logic;
i1 : in  unsigned(0 downto 0);
i2 : in  unsigned(0 downto 0);
i3 : in  unsigned(0 downto 0);
o1 : out unsigned(9 downto 0);
o2 : out unsigned(0 downto 0));
end component cf_fft_2048_16_26;
component cf_fft_2048_16_30 is
port (
clock_c : in std_logic;
i1 : in  unsigned(63 downto 0);
i2 : in  unsigned(0 downto 0);
i3 : in  unsigned(8 downto 0);
i4 : in  unsigned(0 downto 0);
i5 : in  unsigned(0 downto 0);
i6 : in  unsigned(0 downto 0);
o1 : out unsigned(0 downto 0);
o2 : out unsigned(0 downto 0);
o3 : out unsigned(63 downto 0));
end component cf_fft_2048_16_30;
component cf_fft_2048_16_31 is
port (
clock_c : in std_logic;
i1 : in  unsigned(63 downto 0);
i2 : in  unsigned(0 downto 0);
i3 : in  unsigned(8 downto 0);
i4 : in  unsigned(0 downto 0);
i5 : in  unsigned(0 downto 0);
i6 : in  unsigned(0 downto 0);
o1 : out unsigned(63 downto 0));
end component cf_fft_2048_16_31;
begin
n1 <= s27_1(9 downto 9) &
  s27_1(8 downto 8) &
  s27_1(7 downto 7) &
  s27_1(6 downto 6);
n2 <= s26_1 & s26_2;
process (clock_c) begin
  if rising_edge(clock_c) then
    if i5 = "1" then
      n3 <= "0";
    elsif i4 = "1" then
      n3 <= s27_2;
    end if;
  end if;
end process;
process (clock_c) begin
  if rising_edge(clock_c) then
    if i5 = "1" then
      n4 <= "0";
    elsif i4 = "1" then
      n4 <= n3;
    end if;
  end if;
end process;
process (clock_c) begin
  if rising_edge(clock_c) then
    if i5 = "1" then
      n5 <= "0";
    elsif i4 = "1" then
      n5 <= n4;
    end if;
  end if;
end process;
process (clock_c) begin
  if rising_edge(clock_c) then
    if i5 = "1" then
      n6 <= "0";
    elsif i4 = "1" then
      n6 <= n5;
    end if;
  end if;
end process;
n7 <= s27_1(9 downto 9) &
  s27_1(8 downto 8) &
  s27_1(7 downto 7) &
  s27_1(6 downto 6) &
  s27_1(5 downto 5) &
  s27_1(4 downto 4) &
  s27_1(3 downto 3) &
  s27_1(2 downto 2) &
  s27_1(1 downto 1);
process (clock_c) begin
  if rising_edge(clock_c) then
    if i5 = "1" then
      n8 <= "000000000";
    elsif i4 = "1" then
      n8 <= n7;
    end if;
  end if;
end process;
process (clock_c) begin
  if rising_edge(clock_c) then
    if i5 = "1" then
      n9 <= "000000000";
    elsif i4 = "1" then
      n9 <= n8;
    end if;
  end if;
end process;
process (clock_c) begin
  if rising_edge(clock_c) then
    if i5 = "1" then
      n10 <= "000000000";
    elsif i4 = "1" then
      n10 <= n9;
    end if;
  end if;
end process;
process (clock_c) begin
  if rising_edge(clock_c) then
    if i5 = "1" then
      n11 <= "000000000";
    elsif i4 = "1" then
      n11 <= n10;
    end if;
  end if;
end process;
n12 <= s27_1(0 downto 0);
process (clock_c) begin
  if rising_edge(clock_c) then
    if i5 = "1" then
      n13 <= "0";
    elsif i4 = "1" then
      n13 <= n12;
    end if;
  end if;
end process;
process (clock_c) begin
  if rising_edge(clock_c) then
    if i5 = "1" then
      n14 <= "0";
    elsif i4 = "1" then
      n14 <= n13;
    end if;
  end if;
end process;
process (clock_c) begin
  if rising_edge(clock_c) then
    if i5 = "1" then
      n15 <= "0";
    elsif i4 = "1" then
      n15 <= n14;
    end if;
  end if;
end process;
process (clock_c) begin
  if rising_edge(clock_c) then
    if i5 = "1" then
      n16 <= "0";
    elsif i4 = "1" then
      n16 <= n15;
    end if;
  end if;
end process;
n17 <= not n16;
n18 <= s28_2 & s28_1;
n19 <= s28_3(63 downto 63) &
  s28_3(62 downto 62) &
  s28_3(61 downto 61) &
  s28_3(60 downto 60) &
  s28_3(59 downto 59) &
  s28_3(58 downto 58) &
  s28_3(57 downto 57) &
  s28_3(56 downto 56) &
  s28_3(55 downto 55) &
  s28_3(54 downto 54) &
  s28_3(53 downto 53) &
  s28_3(52 downto 52) &
  s28_3(51 downto 51) &
  s28_3(50 downto 50) &
  s28_3(49 downto 49) &
  s28_3(48 downto 48) &
  s28_3(47 downto 47) &
  s28_3(46 downto 46) &
  s28_3(45 downto 45) &
  s28_3(44 downto 44) &
  s28_3(43 downto 43) &
  s28_3(42 downto 42) &
  s28_3(41 downto 41) &
  s28_3(40 downto 40) &
  s28_3(39 downto 39) &
  s28_3(38 downto 38) &
  s28_3(37 downto 37) &
  s28_3(36 downto 36) &
  s28_3(35 downto 35) &
  s28_3(34 downto 34) &
  s28_3(33 downto 33) &
  s28_3(32 downto 32);
n20 <= s28_3(31 downto 31) &
  s28_3(30 downto 30) &
  s28_3(29 downto 29) &
  s28_3(28 downto 28) &
  s28_3(27 downto 27) &
  s28_3(26 downto 26) &
  s28_3(25 downto 25) &
  s28_3(24 downto 24) &
  s28_3(23 downto 23) &
  s28_3(22 downto 22) &
  s28_3(21 downto 21) &
  s28_3(20 downto 20) &
  s28_3(19 downto 19) &
  s28_3(18 downto 18) &
  s28_3(17 downto 17) &
  s28_3(16 downto 16) &
  s28_3(15 downto 15) &
  s28_3(14 downto 14) &
  s28_3(13 downto 13) &
  s28_3(12 downto 12) &
  s28_3(11 downto 11) &
  s28_3(10 downto 10) &
  s28_3(9 downto 9) &
  s28_3(8 downto 8) &
  s28_3(7 downto 7) &
  s28_3(6 downto 6) &
  s28_3(5 downto 5) &
  s28_3(4 downto 4) &
  s28_3(3 downto 3) &
  s28_3(2 downto 2) &
  s28_3(1 downto 1) &
  s28_3(0 downto 0);
n21 <= s29_1(63 downto 63) &
  s29_1(62 downto 62) &
  s29_1(61 downto 61) &
  s29_1(60 downto 60) &
  s29_1(59 downto 59) &
  s29_1(58 downto 58) &
  s29_1(57 downto 57) &
  s29_1(56 downto 56) &
  s29_1(55 downto 55) &
  s29_1(54 downto 54) &
  s29_1(53 downto 53) &
  s29_1(52 downto 52) &
  s29_1(51 downto 51) &
  s29_1(50 downto 50) &
  s29_1(49 downto 49) &
  s29_1(48 downto 48) &
  s29_1(47 downto 47) &
  s29_1(46 downto 46) &
  s29_1(45 downto 45) &
  s29_1(44 downto 44) &
  s29_1(43 downto 43) &
  s29_1(42 downto 42) &
  s29_1(41 downto 41) &
  s29_1(40 downto 40) &
  s29_1(39 downto 39) &
  s29_1(38 downto 38) &
  s29_1(37 downto 37) &
  s29_1(36 downto 36) &
  s29_1(35 downto 35) &
  s29_1(34 downto 34) &
  s29_1(33 downto 33) &
  s29_1(32 downto 32);
n22 <= s29_1(31 downto 31) &
  s29_1(30 downto 30) &
  s29_1(29 downto 29) &
  s29_1(28 downto 28) &
  s29_1(27 downto 27) &
  s29_1(26 downto 26) &
  s29_1(25 downto 25) &
  s29_1(24 downto 24) &
  s29_1(23 downto 23) &
  s29_1(22 downto 22) &
  s29_1(21 downto 21) &
  s29_1(20 downto 20) &
  s29_1(19 downto 19) &
  s29_1(18 downto 18) &
  s29_1(17 downto 17) &
  s29_1(16 downto 16) &
  s29_1(15 downto 15) &
  s29_1(14 downto 14) &
  s29_1(13 downto 13) &
  s29_1(12 downto 12) &
  s29_1(11 downto 11) &
  s29_1(10 downto 10) &
  s29_1(9 downto 9) &
  s29_1(8 downto 8) &
  s29_1(7 downto 7) &
  s29_1(6 downto 6) &
  s29_1(5 downto 5) &
  s29_1(4 downto 4) &
  s29_1(3 downto 3) &
  s29_1(2 downto 2) &
  s29_1(1 downto 1) &
  s29_1(0 downto 0);
n23 <= n20 when s25_1 = "1" else n19;
n24 <= n22 when s25_1 = "1" else n21;
s25 : cf_fft_2048_16_35 port map (clock_c, n18, i4, i5, s25_1);
s26 : cf_fft_2048_16_12 port map (clock_c, i2, i3, n1, i4, i5, s26_1, s26_2);
s27 : cf_fft_2048_16_26 port map (clock_c, i1, i4, i5, s27_1, s27_2);
s28 : cf_fft_2048_16_30 port map (clock_c, n2, n6, n11, n17, i4, i5, s28_1, s28_2, s28_3);
s29 : cf_fft_2048_16_31 port map (clock_c, n2, n6, n11, n16, i4, i5, s29_1);
o3 <= n24;
o2 <= n23;
o1 <= s28_1;
end architecture rtl;

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
entity cf_fft_2048_16_10 is
port (
clock_c : in std_logic;
i1 : in  unsigned(31 downto 0);
i2 : in  unsigned(31 downto 0);
i3 : in  unsigned(2 downto 0);
i4 : in  unsigned(0 downto 0);
i5 : in  unsigned(0 downto 0);
o1 : out unsigned(31 downto 0);
o2 : out unsigned(31 downto 0));
end entity cf_fft_2048_16_10;
architecture rtl of cf_fft_2048_16_10 is
signal n1 : unsigned(31 downto 0) := "00000000000000000000000000000000";
signal n2 : unsigned(15 downto 0);
signal n3 : unsigned(15 downto 0);
signal n4 : unsigned(31 downto 0) := "00000000000000000000000000000000";
signal n5 : unsigned(15 downto 0);
signal n6 : unsigned(15 downto 0);
signal n7 : unsigned(15 downto 0) := "0000000000000000";
signal n8 : unsigned(15 downto 0) := "0000000000000000";
signal n9 : unsigned(15 downto 0) := "0000000000000000";
signal n10 : unsigned(15 downto 0) := "0000000000000000";
signal n11 : unsigned(31 downto 0) := "00000000000000000000000000000000";
signal n12 : unsigned(15 downto 0);
signal n13 : unsigned(15 downto 0);
signal n14 : unsigned(31 downto 0);
signal n15 : unsigned(15 downto 0);
signal n16 : unsigned(15 downto 0) := "0000000000000000";
signal n17 : unsigned(31 downto 0);
signal n18 : unsigned(15 downto 0);
signal n19 : unsigned(15 downto 0) := "0000000000000000";
signal n20 : unsigned(15 downto 0);
signal n21 : unsigned(15 downto 0) := "0000000000000000";
signal n22 : unsigned(31 downto 0);
signal n23 : unsigned(15 downto 0);
signal n24 : unsigned(15 downto 0) := "0000000000000000";
signal n25 : unsigned(31 downto 0);
signal n26 : unsigned(15 downto 0);
signal n27 : unsigned(15 downto 0) := "0000000000000000";
signal n28 : unsigned(15 downto 0);
signal n29 : unsigned(15 downto 0) := "0000000000000000";
signal n30 : unsigned(15 downto 0);
signal n31 : unsigned(15 downto 0);
signal n32 : unsigned(31 downto 0);
signal n33 : unsigned(31 downto 0) := "00000000000000000000000000000000";
signal n34 : unsigned(15 downto 0);
signal n35 : unsigned(15 downto 0);
signal n36 : unsigned(31 downto 0);
signal n37 : unsigned(31 downto 0) := "00000000000000000000000000000000";
begin
process (clock_c) begin
  if rising_edge(clock_c) then
    if i5 = "1" then
      n1 <= "00000000000000000000000000000000";
    elsif i4 = "1" then
      n1 <= i1;
    end if;
  end if;
end process;
n2 <= n1(31 downto 31) &
  n1(30 downto 30) &
  n1(29 downto 29) &
  n1(28 downto 28) &
  n1(27 downto 27) &
  n1(26 downto 26) &
  n1(25 downto 25) &
  n1(24 downto 24) &
  n1(23 downto 23) &
  n1(22 downto 22) &
  n1(21 downto 21) &
  n1(20 downto 20) &
  n1(19 downto 19) &
  n1(18 downto 18) &
  n1(17 downto 17) &
  n1(16 downto 16);
n3 <= n1(15 downto 15) &
  n1(14 downto 14) &
  n1(13 downto 13) &
  n1(12 downto 12) &
  n1(11 downto 11) &
  n1(10 downto 10) &
  n1(9 downto 9) &
  n1(8 downto 8) &
  n1(7 downto 7) &
  n1(6 downto 6) &
  n1(5 downto 5) &
  n1(4 downto 4) &
  n1(3 downto 3) &
  n1(2 downto 2) &
  n1(1 downto 1) &
  n1(0 downto 0);
process (clock_c) begin
  if rising_edge(clock_c) then
    if i5 = "1" then
      n4 <= "00000000000000000000000000000000";
    elsif i4 = "1" then
      n4 <= i2;
    end if;
  end if;
end process;
n5 <= n4(31 downto 31) &
  n4(30 downto 30) &
  n4(29 downto 29) &
  n4(28 downto 28) &
  n4(27 downto 27) &
  n4(26 downto 26) &
  n4(25 downto 25) &
  n4(24 downto 24) &
  n4(23 downto 23) &
  n4(22 downto 22) &
  n4(21 downto 21) &
  n4(20 downto 20) &
  n4(19 downto 19) &
  n4(18 downto 18) &
  n4(17 downto 17) &
  n4(16 downto 16);
n6 <= n4(15 downto 15) &
  n4(14 downto 14) &
  n4(13 downto 13) &
  n4(12 downto 12) &
  n4(11 downto 11) &
  n4(10 downto 10) &
  n4(9 downto 9) &
  n4(8 downto 8) &
  n4(7 downto 7) &
  n4(6 downto 6) &
  n4(5 downto 5) &
  n4(4 downto 4) &
  n4(3 downto 3) &
  n4(2 downto 2) &
  n4(1 downto 1) &
  n4(0 downto 0);
process (clock_c) begin
  if rising_edge(clock_c) then
    if i5 = "1" then
      n7 <= "0000000000000000";
    elsif i4 = "1" then
      n7 <= n2;
    end if;
  end if;
end process;
process (clock_c) begin
  if rising_edge(clock_c) then
    if i5 = "1" then
      n8 <= "0000000000000000";
    elsif i4 = "1" then
      n8 <= n7;
    end if;
  end if;
end process;
process (clock_c) begin
  if rising_edge(clock_c) then
    if i5 = "1" then
      n9 <= "0000000000000000";
    elsif i4 = "1" then
      n9 <= n3;
    end if;
  end if;
end process;
process (clock_c) begin
  if rising_edge(clock_c) then
    if i5 = "1" then
      n10 <= "0000000000000000";
    elsif i4 = "1" then
      n10 <= n9;
    end if;
  end if;
end process;
process (clock_c) begin
  if rising_edge(clock_c) then 
    if i4 = "1" then
      case i3 is
        when "000" => n11 <= "01111111111111110000000000000000";
        when "001" => n11 <= "01110110010000011100111100000100";
        when "010" => n11 <= "01011010100000101010010101111101";
        when "011" => n11 <= "00110000111110111000100110111110";
        when "100" => n11 <= "00000000000000001000000000000000";
        when "101" => n11 <= "11001111000001001000100110111110";
        when "110" => n11 <= "10100101011111011010010101111101";
        when "111" => n11 <= "10001001101111101100111100000100";
        when others => n11 <= "XXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX";
      end case;
    end if;
  end if;
end process;
n12 <= n11(31 downto 31) &
  n11(30 downto 30) &
  n11(29 downto 29) &
  n11(28 downto 28) &
  n11(27 downto 27) &
  n11(26 downto 26) &
  n11(25 downto 25) &
  n11(24 downto 24) &
  n11(23 downto 23) &
  n11(22 downto 22) &
  n11(21 downto 21) &
  n11(20 downto 20) &
  n11(19 downto 19) &
  n11(18 downto 18) &
  n11(17 downto 17) &
  n11(16 downto 16);
n13 <= n11(15 downto 15) &
  n11(14 downto 14) &
  n11(13 downto 13) &
  n11(12 downto 12) &
  n11(11 downto 11) &
  n11(10 downto 10) &
  n11(9 downto 9) &
  n11(8 downto 8) &
  n11(7 downto 7) &
  n11(6 downto 6) &
  n11(5 downto 5) &
  n11(4 downto 4) &
  n11(3 downto 3) &
  n11(2 downto 2) &
  n11(1 downto 1) &
  n11(0 downto 0);
n14 <= unsigned(signed(n5) * signed(n12));
n15 <= n14(30 downto 30) &
  n14(29 downto 29) &
  n14(28 downto 28) &
  n14(27 downto 27) &
  n14(26 downto 26) &
  n14(25 downto 25) &
  n14(24 downto 24) &
  n14(23 downto 23) &
  n14(22 downto 22) &
  n14(21 downto 21) &
  n14(20 downto 20) &
  n14(19 downto 19) &
  n14(18 downto 18) &
  n14(17 downto 17) &
  n14(16 downto 16) &
  n14(15 downto 15);
process (clock_c) begin
  if rising_edge(clock_c) then
    if i5 = "1" then
      n16 <= "0000000000000000";
    elsif i4 = "1" then
      n16 <= n15;
    end if;
  end if;
end process;
n17 <= unsigned(signed(n6) * signed(n13));
n18 <= n17(30 downto 30) &
  n17(29 downto 29) &
  n17(28 downto 28) &
  n17(27 downto 27) &
  n17(26 downto 26) &
  n17(25 downto 25) &
  n17(24 downto 24) &
  n17(23 downto 23) &
  n17(22 downto 22) &
  n17(21 downto 21) &
  n17(20 downto 20) &
  n17(19 downto 19) &
  n17(18 downto 18) &
  n17(17 downto 17) &
  n17(16 downto 16) &
  n17(15 downto 15);
process (clock_c) begin
  if rising_edge(clock_c) then
    if i5 = "1" then
      n19 <= "0000000000000000";
    elsif i4 = "1" then
      n19 <= n18;
    end if;
  end if;
end process;
n20 <= n16 - n19;
process (clock_c) begin
  if rising_edge(clock_c) then
    if i5 = "1" then
      n21 <= "0000000000000000";
    elsif i4 = "1" then
      n21 <= n20;
    end if;
  end if;
end process;
n22 <= unsigned(signed(n5) * signed(n13));
n23 <= n22(30 downto 30) &
  n22(29 downto 29) &
  n22(28 downto 28) &
  n22(27 downto 27) &
  n22(26 downto 26) &
  n22(25 downto 25) &
  n22(24 downto 24) &
  n22(23 downto 23) &
  n22(22 downto 22) &
  n22(21 downto 21) &
  n22(20 downto 20) &
  n22(19 downto 19) &
  n22(18 downto 18) &
  n22(17 downto 17) &
  n22(16 downto 16) &
  n22(15 downto 15);
process (clock_c) begin
  if rising_edge(clock_c) then
    if i5 = "1" then
      n24 <= "0000000000000000";
    elsif i4 = "1" then
      n24 <= n23;
    end if;
  end if;
end process;
n25 <= unsigned(signed(n6) * signed(n12));
n26 <= n25(30 downto 30) &
  n25(29 downto 29) &
  n25(28 downto 28) &
  n25(27 downto 27) &
  n25(26 downto 26) &
  n25(25 downto 25) &
  n25(24 downto 24) &
  n25(23 downto 23) &
  n25(22 downto 22) &
  n25(21 downto 21) &
  n25(20 downto 20) &
  n25(19 downto 19) &
  n25(18 downto 18) &
  n25(17 downto 17) &
  n25(16 downto 16) &
  n25(15 downto 15);
process (clock_c) begin
  if rising_edge(clock_c) then
    if i5 = "1" then
      n27 <= "0000000000000000";
    elsif i4 = "1" then
      n27 <= n26;
    end if;
  end if;
end process;
n28 <= n24 + n27;
process (clock_c) begin
  if rising_edge(clock_c) then
    if i5 = "1" then
      n29 <= "0000000000000000";
    elsif i4 = "1" then
      n29 <= n28;
    end if;
  end if;
end process;
n30 <= n8 + n21;
n31 <= n10 + n29;
n32 <= n30 & n31;
process (clock_c) begin
  if rising_edge(clock_c) then
    if i5 = "1" then
      n33 <= "00000000000000000000000000000000";
    elsif i4 = "1" then
      n33 <= n32;
    end if;
  end if;
end process;
n34 <= n8 - n21;
n35 <= n10 - n29;
n36 <= n34 & n35;
process (clock_c) begin
  if rising_edge(clock_c) then
    if i5 = "1" then
      n37 <= "00000000000000000000000000000000";
    elsif i4 = "1" then
      n37 <= n36;
    end if;
  end if;
end process;
o2 <= n37;
o1 <= n33;
end architecture rtl;

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
entity cf_fft_2048_16_9 is
port (
clock_c : in std_logic;
i1 : in  unsigned(0 downto 0);
i2 : in  unsigned(31 downto 0);
i3 : in  unsigned(31 downto 0);
i4 : in  unsigned(0 downto 0);
i5 : in  unsigned(0 downto 0);
o1 : out unsigned(0 downto 0);
o2 : out unsigned(31 downto 0);
o3 : out unsigned(31 downto 0));
end entity cf_fft_2048_16_9;
architecture rtl of cf_fft_2048_16_9 is
signal n1 : unsigned(2 downto 0);
signal n2 : unsigned(63 downto 0);
signal n3 : unsigned(0 downto 0) := "0";
signal n4 : unsigned(0 downto 0) := "0";
signal n5 : unsigned(0 downto 0) := "0";
signal n6 : unsigned(0 downto 0) := "0";
signal n7 : unsigned(8 downto 0);
signal n8 : unsigned(8 downto 0) := "000000000";
signal n9 : unsigned(8 downto 0) := "000000000";
signal n10 : unsigned(8 downto 0) := "000000000";
signal n11 : unsigned(8 downto 0) := "000000000";
signal n12 : unsigned(0 downto 0);
signal n13 : unsigned(0 downto 0) := "0";
signal n14 : unsigned(0 downto 0) := "0";
signal n15 : unsigned(0 downto 0) := "0";
signal n16 : unsigned(0 downto 0) := "0";
signal n17 : unsigned(0 downto 0);
signal n18 : unsigned(1 downto 0);
signal n19 : unsigned(31 downto 0);
signal n20 : unsigned(31 downto 0);
signal n21 : unsigned(31 downto 0);
signal n22 : unsigned(31 downto 0);
signal n23 : unsigned(31 downto 0);
signal n24 : unsigned(31 downto 0);
signal s25_1 : unsigned(31 downto 0);
signal s25_2 : unsigned(31 downto 0);
signal s26_1 : unsigned(0 downto 0);
signal s27_1 : unsigned(0 downto 0);
signal s27_2 : unsigned(0 downto 0);
signal s27_3 : unsigned(63 downto 0);
signal s28_1 : unsigned(63 downto 0);
signal s29_1 : unsigned(9 downto 0);
signal s29_2 : unsigned(0 downto 0);
component cf_fft_2048_16_10 is
port (
clock_c : in std_logic;
i1 : in  unsigned(31 downto 0);
i2 : in  unsigned(31 downto 0);
i3 : in  unsigned(2 downto 0);
i4 : in  unsigned(0 downto 0);
i5 : in  unsigned(0 downto 0);
o1 : out unsigned(31 downto 0);
o2 : out unsigned(31 downto 0));
end component cf_fft_2048_16_10;
component cf_fft_2048_16_35 is
port (
clock_c : in std_logic;
i1 : in  unsigned(1 downto 0);
i2 : in  unsigned(0 downto 0);
i3 : in  unsigned(0 downto 0);
o1 : out unsigned(0 downto 0));
end component cf_fft_2048_16_35;
component cf_fft_2048_16_30 is
port (
clock_c : in std_logic;
i1 : in  unsigned(63 downto 0);
i2 : in  unsigned(0 downto 0);
i3 : in  unsigned(8 downto 0);
i4 : in  unsigned(0 downto 0);
i5 : in  unsigned(0 downto 0);
i6 : in  unsigned(0 downto 0);
o1 : out unsigned(0 downto 0);
o2 : out unsigned(0 downto 0);
o3 : out unsigned(63 downto 0));
end component cf_fft_2048_16_30;
component cf_fft_2048_16_31 is
port (
clock_c : in std_logic;
i1 : in  unsigned(63 downto 0);
i2 : in  unsigned(0 downto 0);
i3 : in  unsigned(8 downto 0);
i4 : in  unsigned(0 downto 0);
i5 : in  unsigned(0 downto 0);
i6 : in  unsigned(0 downto 0);
o1 : out unsigned(63 downto 0));
end component cf_fft_2048_16_31;
component cf_fft_2048_16_26 is
port (
clock_c : in std_logic;
i1 : in  unsigned(0 downto 0);
i2 : in  unsigned(0 downto 0);
i3 : in  unsigned(0 downto 0);
o1 : out unsigned(9 downto 0);
o2 : out unsigned(0 downto 0));
end component cf_fft_2048_16_26;
begin
n1 <= s29_1(9 downto 9) &
  s29_1(8 downto 8) &
  s29_1(7 downto 7);
n2 <= s25_1 & s25_2;
process (clock_c) begin
  if rising_edge(clock_c) then
    if i5 = "1" then
      n3 <= "0";
    elsif i4 = "1" then
      n3 <= s29_2;
    end if;
  end if;
end process;
process (clock_c) begin
  if rising_edge(clock_c) then
    if i5 = "1" then
      n4 <= "0";
    elsif i4 = "1" then
      n4 <= n3;
    end if;
  end if;
end process;
process (clock_c) begin
  if rising_edge(clock_c) then
    if i5 = "1" then
      n5 <= "0";
    elsif i4 = "1" then
      n5 <= n4;
    end if;
  end if;
end process;
process (clock_c) begin
  if rising_edge(clock_c) then
    if i5 = "1" then
      n6 <= "0";
    elsif i4 = "1" then
      n6 <= n5;
    end if;
  end if;
end process;
n7 <= s29_1(9 downto 9) &
  s29_1(8 downto 8) &
  s29_1(7 downto 7) &
  s29_1(6 downto 6) &
  s29_1(5 downto 5) &
  s29_1(4 downto 4) &
  s29_1(3 downto 3) &
  s29_1(2 downto 2) &
  s29_1(1 downto 1);
process (clock_c) begin
  if rising_edge(clock_c) then
    if i5 = "1" then
      n8 <= "000000000";
    elsif i4 = "1" then
      n8 <= n7;
    end if;
  end if;
end process;
process (clock_c) begin
  if rising_edge(clock_c) then
    if i5 = "1" then
      n9 <= "000000000";
    elsif i4 = "1" then
      n9 <= n8;
    end if;
  end if;
end process;
process (clock_c) begin
  if rising_edge(clock_c) then
    if i5 = "1" then
      n10 <= "000000000";
    elsif i4 = "1" then
      n10 <= n9;
    end if;
  end if;
end process;
process (clock_c) begin
  if rising_edge(clock_c) then
    if i5 = "1" then
      n11 <= "000000000";
    elsif i4 = "1" then
      n11 <= n10;
    end if;
  end if;
end process;
n12 <= s29_1(0 downto 0);
process (clock_c) begin
  if rising_edge(clock_c) then
    if i5 = "1" then
      n13 <= "0";
    elsif i4 = "1" then
      n13 <= n12;
    end if;
  end if;
end process;
process (clock_c) begin
  if rising_edge(clock_c) then
    if i5 = "1" then
      n14 <= "0";
    elsif i4 = "1" then
      n14 <= n13;
    end if;
  end if;
end process;
process (clock_c) begin
  if rising_edge(clock_c) then
    if i5 = "1" then
      n15 <= "0";
    elsif i4 = "1" then
      n15 <= n14;
    end if;
  end if;
end process;
process (clock_c) begin
  if rising_edge(clock_c) then
    if i5 = "1" then
      n16 <= "0";
    elsif i4 = "1" then
      n16 <= n15;
    end if;
  end if;
end process;
n17 <= not n16;
n18 <= s27_2 & s27_1;
n19 <= s27_3(63 downto 63) &
  s27_3(62 downto 62) &
  s27_3(61 downto 61) &
  s27_3(60 downto 60) &
  s27_3(59 downto 59) &
  s27_3(58 downto 58) &
  s27_3(57 downto 57) &
  s27_3(56 downto 56) &
  s27_3(55 downto 55) &
  s27_3(54 downto 54) &
  s27_3(53 downto 53) &
  s27_3(52 downto 52) &
  s27_3(51 downto 51) &
  s27_3(50 downto 50) &
  s27_3(49 downto 49) &
  s27_3(48 downto 48) &
  s27_3(47 downto 47) &
  s27_3(46 downto 46) &
  s27_3(45 downto 45) &
  s27_3(44 downto 44) &
  s27_3(43 downto 43) &
  s27_3(42 downto 42) &
  s27_3(41 downto 41) &
  s27_3(40 downto 40) &
  s27_3(39 downto 39) &
  s27_3(38 downto 38) &
  s27_3(37 downto 37) &
  s27_3(36 downto 36) &
  s27_3(35 downto 35) &
  s27_3(34 downto 34) &
  s27_3(33 downto 33) &
  s27_3(32 downto 32);
n20 <= s27_3(31 downto 31) &
  s27_3(30 downto 30) &
  s27_3(29 downto 29) &
  s27_3(28 downto 28) &
  s27_3(27 downto 27) &
  s27_3(26 downto 26) &
  s27_3(25 downto 25) &
  s27_3(24 downto 24) &
  s27_3(23 downto 23) &
  s27_3(22 downto 22) &
  s27_3(21 downto 21) &
  s27_3(20 downto 20) &
  s27_3(19 downto 19) &
  s27_3(18 downto 18) &
  s27_3(17 downto 17) &
  s27_3(16 downto 16) &
  s27_3(15 downto 15) &
  s27_3(14 downto 14) &
  s27_3(13 downto 13) &
  s27_3(12 downto 12) &
  s27_3(11 downto 11) &
  s27_3(10 downto 10) &
  s27_3(9 downto 9) &
  s27_3(8 downto 8) &
  s27_3(7 downto 7) &
  s27_3(6 downto 6) &
  s27_3(5 downto 5) &
  s27_3(4 downto 4) &
  s27_3(3 downto 3) &
  s27_3(2 downto 2) &
  s27_3(1 downto 1) &
  s27_3(0 downto 0);
n21 <= s28_1(63 downto 63) &
  s28_1(62 downto 62) &
  s28_1(61 downto 61) &
  s28_1(60 downto 60) &
  s28_1(59 downto 59) &
  s28_1(58 downto 58) &
  s28_1(57 downto 57) &
  s28_1(56 downto 56) &
  s28_1(55 downto 55) &
  s28_1(54 downto 54) &
  s28_1(53 downto 53) &
  s28_1(52 downto 52) &
  s28_1(51 downto 51) &
  s28_1(50 downto 50) &
  s28_1(49 downto 49) &
  s28_1(48 downto 48) &
  s28_1(47 downto 47) &
  s28_1(46 downto 46) &
  s28_1(45 downto 45) &
  s28_1(44 downto 44) &
  s28_1(43 downto 43) &
  s28_1(42 downto 42) &
  s28_1(41 downto 41) &
  s28_1(40 downto 40) &
  s28_1(39 downto 39) &
  s28_1(38 downto 38) &
  s28_1(37 downto 37) &
  s28_1(36 downto 36) &
  s28_1(35 downto 35) &
  s28_1(34 downto 34) &
  s28_1(33 downto 33) &
  s28_1(32 downto 32);
n22 <= s28_1(31 downto 31) &
  s28_1(30 downto 30) &
  s28_1(29 downto 29) &
  s28_1(28 downto 28) &
  s28_1(27 downto 27) &
  s28_1(26 downto 26) &
  s28_1(25 downto 25) &
  s28_1(24 downto 24) &
  s28_1(23 downto 23) &
  s28_1(22 downto 22) &
  s28_1(21 downto 21) &
  s28_1(20 downto 20) &
  s28_1(19 downto 19) &
  s28_1(18 downto 18) &
  s28_1(17 downto 17) &
  s28_1(16 downto 16) &
  s28_1(15 downto 15) &
  s28_1(14 downto 14) &
  s28_1(13 downto 13) &
  s28_1(12 downto 12) &
  s28_1(11 downto 11) &
  s28_1(10 downto 10) &
  s28_1(9 downto 9) &
  s28_1(8 downto 8) &
  s28_1(7 downto 7) &
  s28_1(6 downto 6) &
  s28_1(5 downto 5) &
  s28_1(4 downto 4) &
  s28_1(3 downto 3) &
  s28_1(2 downto 2) &
  s28_1(1 downto 1) &
  s28_1(0 downto 0);
n23 <= n20 when s26_1 = "1" else n19;
n24 <= n22 when s26_1 = "1" else n21;
s25 : cf_fft_2048_16_10 port map (clock_c, i2, i3, n1, i4, i5, s25_1, s25_2);
s26 : cf_fft_2048_16_35 port map (clock_c, n18, i4, i5, s26_1);
s27 : cf_fft_2048_16_30 port map (clock_c, n2, n6, n11, n17, i4, i5, s27_1, s27_2, s27_3);
s28 : cf_fft_2048_16_31 port map (clock_c, n2, n6, n11, n16, i4, i5, s28_1);
s29 : cf_fft_2048_16_26 port map (clock_c, i1, i4, i5, s29_1, s29_2);
o3 <= n24;
o2 <= n23;
o1 <= s27_1;
end architecture rtl;

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
entity cf_fft_2048_16_8 is
port (
clock_c : in std_logic;
i1 : in  unsigned(0 downto 0);
i2 : in  unsigned(31 downto 0);
i3 : in  unsigned(31 downto 0);
i4 : in  unsigned(0 downto 0);
i5 : in  unsigned(0 downto 0);
o1 : out unsigned(0 downto 0);
o2 : out unsigned(31 downto 0);
o3 : out unsigned(31 downto 0));
end entity cf_fft_2048_16_8;
architecture rtl of cf_fft_2048_16_8 is
signal s1_1 : unsigned(0 downto 0);
signal s1_2 : unsigned(31 downto 0);
signal s1_3 : unsigned(31 downto 0);
signal s2_1 : unsigned(0 downto 0);
signal s2_2 : unsigned(31 downto 0);
signal s2_3 : unsigned(31 downto 0);
signal s3_1 : unsigned(0 downto 0);
signal s3_2 : unsigned(31 downto 0);
signal s3_3 : unsigned(31 downto 0);
signal s4_1 : unsigned(0 downto 0);
signal s4_2 : unsigned(31 downto 0);
signal s4_3 : unsigned(31 downto 0);
signal s5_1 : unsigned(0 downto 0);
signal s5_2 : unsigned(31 downto 0);
signal s5_3 : unsigned(31 downto 0);
signal s6_1 : unsigned(0 downto 0);
signal s6_2 : unsigned(31 downto 0);
signal s6_3 : unsigned(31 downto 0);
signal s7_1 : unsigned(0 downto 0);
signal s7_2 : unsigned(31 downto 0);
signal s7_3 : unsigned(31 downto 0);
signal s8_1 : unsigned(0 downto 0);
signal s8_2 : unsigned(31 downto 0);
signal s8_3 : unsigned(31 downto 0);
component cf_fft_2048_16_23 is
port (
clock_c : in std_logic;
i1 : in  unsigned(0 downto 0);
i2 : in  unsigned(31 downto 0);
i3 : in  unsigned(31 downto 0);
i4 : in  unsigned(0 downto 0);
i5 : in  unsigned(0 downto 0);
o1 : out unsigned(0 downto 0);
o2 : out unsigned(31 downto 0);
o3 : out unsigned(31 downto 0));
end component cf_fft_2048_16_23;
component cf_fft_2048_16_21 is
port (
clock_c : in std_logic;
i1 : in  unsigned(0 downto 0);
i2 : in  unsigned(31 downto 0);
i3 : in  unsigned(31 downto 0);
i4 : in  unsigned(0 downto 0);
i5 : in  unsigned(0 downto 0);
o1 : out unsigned(0 downto 0);
o2 : out unsigned(31 downto 0);
o3 : out unsigned(31 downto 0));
end component cf_fft_2048_16_21;
component cf_fft_2048_16_19 is
port (
clock_c : in std_logic;
i1 : in  unsigned(0 downto 0);
i2 : in  unsigned(31 downto 0);
i3 : in  unsigned(31 downto 0);
i4 : in  unsigned(0 downto 0);
i5 : in  unsigned(0 downto 0);
o1 : out unsigned(0 downto 0);
o2 : out unsigned(31 downto 0);
o3 : out unsigned(31 downto 0));
end component cf_fft_2048_16_19;
component cf_fft_2048_16_17 is
port (
clock_c : in std_logic;
i1 : in  unsigned(0 downto 0);
i2 : in  unsigned(31 downto 0);
i3 : in  unsigned(31 downto 0);
i4 : in  unsigned(0 downto 0);
i5 : in  unsigned(0 downto 0);
o1 : out unsigned(0 downto 0);
o2 : out unsigned(31 downto 0);
o3 : out unsigned(31 downto 0));
end component cf_fft_2048_16_17;
component cf_fft_2048_16_15 is
port (
clock_c : in std_logic;
i1 : in  unsigned(0 downto 0);
i2 : in  unsigned(31 downto 0);
i3 : in  unsigned(31 downto 0);
i4 : in  unsigned(0 downto 0);
i5 : in  unsigned(0 downto 0);
o1 : out unsigned(0 downto 0);
o2 : out unsigned(31 downto 0);
o3 : out unsigned(31 downto 0));
end component cf_fft_2048_16_15;
component cf_fft_2048_16_13 is
port (
clock_c : in std_logic;
i1 : in  unsigned(0 downto 0);
i2 : in  unsigned(31 downto 0);
i3 : in  unsigned(31 downto 0);
i4 : in  unsigned(0 downto 0);
i5 : in  unsigned(0 downto 0);
o1 : out unsigned(0 downto 0);
o2 : out unsigned(31 downto 0);
o3 : out unsigned(31 downto 0));
end component cf_fft_2048_16_13;
component cf_fft_2048_16_11 is
port (
clock_c : in std_logic;
i1 : in  unsigned(0 downto 0);
i2 : in  unsigned(31 downto 0);
i3 : in  unsigned(31 downto 0);
i4 : in  unsigned(0 downto 0);
i5 : in  unsigned(0 downto 0);
o1 : out unsigned(0 downto 0);
o2 : out unsigned(31 downto 0);
o3 : out unsigned(31 downto 0));
end component cf_fft_2048_16_11;
component cf_fft_2048_16_9 is
port (
clock_c : in std_logic;
i1 : in  unsigned(0 downto 0);
i2 : in  unsigned(31 downto 0);
i3 : in  unsigned(31 downto 0);
i4 : in  unsigned(0 downto 0);
i5 : in  unsigned(0 downto 0);
o1 : out unsigned(0 downto 0);
o2 : out unsigned(31 downto 0);
o3 : out unsigned(31 downto 0));
end component cf_fft_2048_16_9;
begin
s1 : cf_fft_2048_16_23 port map (clock_c, s2_1, s2_2, s2_3, i4, i5, s1_1, s1_2, s1_3);
s2 : cf_fft_2048_16_21 port map (clock_c, s3_1, s3_2, s3_3, i4, i5, s2_1, s2_2, s2_3);
s3 : cf_fft_2048_16_19 port map (clock_c, s4_1, s4_2, s4_3, i4, i5, s3_1, s3_2, s3_3);
s4 : cf_fft_2048_16_17 port map (clock_c, s5_1, s5_2, s5_3, i4, i5, s4_1, s4_2, s4_3);
s5 : cf_fft_2048_16_15 port map (clock_c, s6_1, s6_2, s6_3, i4, i5, s5_1, s5_2, s5_3);
s6 : cf_fft_2048_16_13 port map (clock_c, s7_1, s7_2, s7_3, i4, i5, s6_1, s6_2, s6_3);
s7 : cf_fft_2048_16_11 port map (clock_c, s8_1, s8_2, s8_3, i4, i5, s7_1, s7_2, s7_3);
s8 : cf_fft_2048_16_9 port map (clock_c, i1, i2, i3, i4, i5, s8_1, s8_2, s8_3);
o3 <= s1_3;
o2 <= s1_2;
o1 <= s1_1;
end architecture rtl;

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
entity cf_fft_2048_16_7 is
port (
clock_c : in std_logic;
i1 : in  unsigned(31 downto 0);
i2 : in  unsigned(31 downto 0);
i3 : in  unsigned(0 downto 0);
i4 : in  unsigned(0 downto 0);
i5 : in  unsigned(0 downto 0);
o1 : out unsigned(31 downto 0);
o2 : out unsigned(31 downto 0));
end entity cf_fft_2048_16_7;
architecture rtl of cf_fft_2048_16_7 is
signal n1 : unsigned(31 downto 0) := "00000000000000000000000000000000";
signal n2 : unsigned(15 downto 0);
signal n3 : unsigned(15 downto 0);
signal n4 : unsigned(31 downto 0) := "00000000000000000000000000000000";
signal n5 : unsigned(15 downto 0);
signal n6 : unsigned(15 downto 0);
signal n7 : unsigned(15 downto 0) := "0000000000000000";
signal n8 : unsigned(15 downto 0) := "0000000000000000";
signal n9 : unsigned(15 downto 0) := "0000000000000000";
signal n10 : unsigned(15 downto 0) := "0000000000000000";
signal n11 : unsigned(31 downto 0) := "00000000000000000000000000000000";
signal n12 : unsigned(15 downto 0);
signal n13 : unsigned(15 downto 0);
signal n14 : unsigned(31 downto 0);
signal n15 : unsigned(15 downto 0);
signal n16 : unsigned(15 downto 0) := "0000000000000000";
signal n17 : unsigned(31 downto 0);
signal n18 : unsigned(15 downto 0);
signal n19 : unsigned(15 downto 0) := "0000000000000000";
signal n20 : unsigned(15 downto 0);
signal n21 : unsigned(15 downto 0) := "0000000000000000";
signal n22 : unsigned(31 downto 0);
signal n23 : unsigned(15 downto 0);
signal n24 : unsigned(15 downto 0) := "0000000000000000";
signal n25 : unsigned(31 downto 0);
signal n26 : unsigned(15 downto 0);
signal n27 : unsigned(15 downto 0) := "0000000000000000";
signal n28 : unsigned(15 downto 0);
signal n29 : unsigned(15 downto 0) := "0000000000000000";
signal n30 : unsigned(15 downto 0);
signal n31 : unsigned(15 downto 0);
signal n32 : unsigned(31 downto 0);
signal n33 : unsigned(31 downto 0) := "00000000000000000000000000000000";
signal n34 : unsigned(15 downto 0);
signal n35 : unsigned(15 downto 0);
signal n36 : unsigned(31 downto 0);
signal n37 : unsigned(31 downto 0) := "00000000000000000000000000000000";
begin
process (clock_c) begin
  if rising_edge(clock_c) then
    if i5 = "1" then
      n1 <= "00000000000000000000000000000000";
    elsif i4 = "1" then
      n1 <= i1;
    end if;
  end if;
end process;
n2 <= n1(31 downto 31) &
  n1(30 downto 30) &
  n1(29 downto 29) &
  n1(28 downto 28) &
  n1(27 downto 27) &
  n1(26 downto 26) &
  n1(25 downto 25) &
  n1(24 downto 24) &
  n1(23 downto 23) &
  n1(22 downto 22) &
  n1(21 downto 21) &
  n1(20 downto 20) &
  n1(19 downto 19) &
  n1(18 downto 18) &
  n1(17 downto 17) &
  n1(16 downto 16);
n3 <= n1(15 downto 15) &
  n1(14 downto 14) &
  n1(13 downto 13) &
  n1(12 downto 12) &
  n1(11 downto 11) &
  n1(10 downto 10) &
  n1(9 downto 9) &
  n1(8 downto 8) &
  n1(7 downto 7) &
  n1(6 downto 6) &
  n1(5 downto 5) &
  n1(4 downto 4) &
  n1(3 downto 3) &
  n1(2 downto 2) &
  n1(1 downto 1) &
  n1(0 downto 0);
process (clock_c) begin
  if rising_edge(clock_c) then
    if i5 = "1" then
      n4 <= "00000000000000000000000000000000";
    elsif i4 = "1" then
      n4 <= i2;
    end if;
  end if;
end process;
n5 <= n4(31 downto 31) &
  n4(30 downto 30) &
  n4(29 downto 29) &
  n4(28 downto 28) &
  n4(27 downto 27) &
  n4(26 downto 26) &
  n4(25 downto 25) &
  n4(24 downto 24) &
  n4(23 downto 23) &
  n4(22 downto 22) &
  n4(21 downto 21) &
  n4(20 downto 20) &
  n4(19 downto 19) &
  n4(18 downto 18) &
  n4(17 downto 17) &
  n4(16 downto 16);
n6 <= n4(15 downto 15) &
  n4(14 downto 14) &
  n4(13 downto 13) &
  n4(12 downto 12) &
  n4(11 downto 11) &
  n4(10 downto 10) &
  n4(9 downto 9) &
  n4(8 downto 8) &
  n4(7 downto 7) &
  n4(6 downto 6) &
  n4(5 downto 5) &
  n4(4 downto 4) &
  n4(3 downto 3) &
  n4(2 downto 2) &
  n4(1 downto 1) &
  n4(0 downto 0);
process (clock_c) begin
  if rising_edge(clock_c) then
    if i5 = "1" then
      n7 <= "0000000000000000";
    elsif i4 = "1" then
      n7 <= n2;
    end if;
  end if;
end process;
process (clock_c) begin
  if rising_edge(clock_c) then
    if i5 = "1" then
      n8 <= "0000000000000000";
    elsif i4 = "1" then
      n8 <= n7;
    end if;
  end if;
end process;
process (clock_c) begin
  if rising_edge(clock_c) then
    if i5 = "1" then
      n9 <= "0000000000000000";
    elsif i4 = "1" then
      n9 <= n3;
    end if;
  end if;
end process;
process (clock_c) begin
  if rising_edge(clock_c) then
    if i5 = "1" then
      n10 <= "0000000000000000";
    elsif i4 = "1" then
      n10 <= n9;
    end if;
  end if;
end process;
process (clock_c) begin
  if rising_edge(clock_c) then 
    if i4 = "1" then
      case i3 is
        when "0" => n11 <= "01111111111111110000000000000000";
        when "1" => n11 <= "00000000000000001000000000000000";
        when others => n11 <= "XXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX";
      end case;
    end if;
  end if;
end process;
n12 <= n11(31 downto 31) &
  n11(30 downto 30) &
  n11(29 downto 29) &
  n11(28 downto 28) &
  n11(27 downto 27) &
  n11(26 downto 26) &
  n11(25 downto 25) &
  n11(24 downto 24) &
  n11(23 downto 23) &
  n11(22 downto 22) &
  n11(21 downto 21) &
  n11(20 downto 20) &
  n11(19 downto 19) &
  n11(18 downto 18) &
  n11(17 downto 17) &
  n11(16 downto 16);
n13 <= n11(15 downto 15) &
  n11(14 downto 14) &
  n11(13 downto 13) &
  n11(12 downto 12) &
  n11(11 downto 11) &
  n11(10 downto 10) &
  n11(9 downto 9) &
  n11(8 downto 8) &
  n11(7 downto 7) &
  n11(6 downto 6) &
  n11(5 downto 5) &
  n11(4 downto 4) &
  n11(3 downto 3) &
  n11(2 downto 2) &
  n11(1 downto 1) &
  n11(0 downto 0);
n14 <= unsigned(signed(n5) * signed(n12));
n15 <= n14(30 downto 30) &
  n14(29 downto 29) &
  n14(28 downto 28) &
  n14(27 downto 27) &
  n14(26 downto 26) &
  n14(25 downto 25) &
  n14(24 downto 24) &
  n14(23 downto 23) &
  n14(22 downto 22) &
  n14(21 downto 21) &
  n14(20 downto 20) &
  n14(19 downto 19) &
  n14(18 downto 18) &
  n14(17 downto 17) &
  n14(16 downto 16) &
  n14(15 downto 15);
process (clock_c) begin
  if rising_edge(clock_c) then
    if i5 = "1" then
      n16 <= "0000000000000000";
    elsif i4 = "1" then
      n16 <= n15;
    end if;
  end if;
end process;
n17 <= unsigned(signed(n6) * signed(n13));
n18 <= n17(30 downto 30) &
  n17(29 downto 29) &
  n17(28 downto 28) &
  n17(27 downto 27) &
  n17(26 downto 26) &
  n17(25 downto 25) &
  n17(24 downto 24) &
  n17(23 downto 23) &
  n17(22 downto 22) &
  n17(21 downto 21) &
  n17(20 downto 20) &
  n17(19 downto 19) &
  n17(18 downto 18) &
  n17(17 downto 17) &
  n17(16 downto 16) &
  n17(15 downto 15);
process (clock_c) begin
  if rising_edge(clock_c) then
    if i5 = "1" then
      n19 <= "0000000000000000";
    elsif i4 = "1" then
      n19 <= n18;
    end if;
  end if;
end process;
n20 <= n16 - n19;
process (clock_c) begin
  if rising_edge(clock_c) then
    if i5 = "1" then
      n21 <= "0000000000000000";
    elsif i4 = "1" then
      n21 <= n20;
    end if;
  end if;
end process;
n22 <= unsigned(signed(n5) * signed(n13));
n23 <= n22(30 downto 30) &
  n22(29 downto 29) &
  n22(28 downto 28) &
  n22(27 downto 27) &
  n22(26 downto 26) &
  n22(25 downto 25) &
  n22(24 downto 24) &
  n22(23 downto 23) &
  n22(22 downto 22) &
  n22(21 downto 21) &
  n22(20 downto 20) &
  n22(19 downto 19) &
  n22(18 downto 18) &
  n22(17 downto 17) &
  n22(16 downto 16) &
  n22(15 downto 15);
process (clock_c) begin
  if rising_edge(clock_c) then
    if i5 = "1" then
      n24 <= "0000000000000000";
    elsif i4 = "1" then
      n24 <= n23;
    end if;
  end if;
end process;
n25 <= unsigned(signed(n6) * signed(n12));
n26 <= n25(30 downto 30) &
  n25(29 downto 29) &
  n25(28 downto 28) &
  n25(27 downto 27) &
  n25(26 downto 26) &
  n25(25 downto 25) &
  n25(24 downto 24) &
  n25(23 downto 23) &
  n25(22 downto 22) &
  n25(21 downto 21) &
  n25(20 downto 20) &
  n25(19 downto 19) &
  n25(18 downto 18) &
  n25(17 downto 17) &
  n25(16 downto 16) &
  n25(15 downto 15);
process (clock_c) begin
  if rising_edge(clock_c) then
    if i5 = "1" then
      n27 <= "0000000000000000";
    elsif i4 = "1" then
      n27 <= n26;
    end if;
  end if;
end process;
n28 <= n24 + n27;
process (clock_c) begin
  if rising_edge(clock_c) then
    if i5 = "1" then
      n29 <= "0000000000000000";
    elsif i4 = "1" then
      n29 <= n28;
    end if;
  end if;
end process;
n30 <= n8 + n21;
n31 <= n10 + n29;
n32 <= n30 & n31;
process (clock_c) begin
  if rising_edge(clock_c) then
    if i5 = "1" then
      n33 <= "00000000000000000000000000000000";
    elsif i4 = "1" then
      n33 <= n32;
    end if;
  end if;
end process;
n34 <= n8 - n21;
n35 <= n10 - n29;
n36 <= n34 & n35;
process (clock_c) begin
  if rising_edge(clock_c) then
    if i5 = "1" then
      n37 <= "00000000000000000000000000000000";
    elsif i4 = "1" then
      n37 <= n36;
    end if;
  end if;
end process;
o2 <= n37;
o1 <= n33;
end architecture rtl;

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
entity cf_fft_2048_16_6 is
port (
clock_c : in std_logic;
i1 : in  unsigned(0 downto 0);
i2 : in  unsigned(31 downto 0);
i3 : in  unsigned(31 downto 0);
i4 : in  unsigned(0 downto 0);
i5 : in  unsigned(0 downto 0);
o1 : out unsigned(0 downto 0);
o2 : out unsigned(31 downto 0);
o3 : out unsigned(31 downto 0));
end entity cf_fft_2048_16_6;
architecture rtl of cf_fft_2048_16_6 is
signal n1 : unsigned(0 downto 0);
signal n2 : unsigned(63 downto 0);
signal n3 : unsigned(0 downto 0) := "0";
signal n4 : unsigned(0 downto 0) := "0";
signal n5 : unsigned(0 downto 0) := "0";
signal n6 : unsigned(0 downto 0) := "0";
signal n7 : unsigned(8 downto 0);
signal n8 : unsigned(8 downto 0) := "000000000";
signal n9 : unsigned(8 downto 0) := "000000000";
signal n10 : unsigned(8 downto 0) := "000000000";
signal n11 : unsigned(8 downto 0) := "000000000";
signal n12 : unsigned(0 downto 0);
signal n13 : unsigned(0 downto 0) := "0";
signal n14 : unsigned(0 downto 0) := "0";
signal n15 : unsigned(0 downto 0) := "0";
signal n16 : unsigned(0 downto 0) := "0";
signal n17 : unsigned(0 downto 0);
signal n18 : unsigned(1 downto 0);
signal n19 : unsigned(31 downto 0);
signal n20 : unsigned(31 downto 0);
signal n21 : unsigned(31 downto 0);
signal n22 : unsigned(31 downto 0);
signal n23 : unsigned(31 downto 0);
signal n24 : unsigned(31 downto 0);
signal s25_1 : unsigned(31 downto 0);
signal s25_2 : unsigned(31 downto 0);
signal s26_1 : unsigned(0 downto 0);
signal s27_1 : unsigned(63 downto 0);
signal s28_1 : unsigned(0 downto 0);
signal s28_2 : unsigned(0 downto 0);
signal s28_3 : unsigned(63 downto 0);
signal s29_1 : unsigned(9 downto 0);
signal s29_2 : unsigned(0 downto 0);
component cf_fft_2048_16_7 is
port (
clock_c : in std_logic;
i1 : in  unsigned(31 downto 0);
i2 : in  unsigned(31 downto 0);
i3 : in  unsigned(0 downto 0);
i4 : in  unsigned(0 downto 0);
i5 : in  unsigned(0 downto 0);
o1 : out unsigned(31 downto 0);
o2 : out unsigned(31 downto 0));
end component cf_fft_2048_16_7;
component cf_fft_2048_16_35 is
port (
clock_c : in std_logic;
i1 : in  unsigned(1 downto 0);
i2 : in  unsigned(0 downto 0);
i3 : in  unsigned(0 downto 0);
o1 : out unsigned(0 downto 0));
end component cf_fft_2048_16_35;
component cf_fft_2048_16_31 is
port (
clock_c : in std_logic;
i1 : in  unsigned(63 downto 0);
i2 : in  unsigned(0 downto 0);
i3 : in  unsigned(8 downto 0);
i4 : in  unsigned(0 downto 0);
i5 : in  unsigned(0 downto 0);
i6 : in  unsigned(0 downto 0);
o1 : out unsigned(63 downto 0));
end component cf_fft_2048_16_31;
component cf_fft_2048_16_30 is
port (
clock_c : in std_logic;
i1 : in  unsigned(63 downto 0);
i2 : in  unsigned(0 downto 0);
i3 : in  unsigned(8 downto 0);
i4 : in  unsigned(0 downto 0);
i5 : in  unsigned(0 downto 0);
i6 : in  unsigned(0 downto 0);
o1 : out unsigned(0 downto 0);
o2 : out unsigned(0 downto 0);
o3 : out unsigned(63 downto 0));
end component cf_fft_2048_16_30;
component cf_fft_2048_16_26 is
port (
clock_c : in std_logic;
i1 : in  unsigned(0 downto 0);
i2 : in  unsigned(0 downto 0);
i3 : in  unsigned(0 downto 0);
o1 : out unsigned(9 downto 0);
o2 : out unsigned(0 downto 0));
end component cf_fft_2048_16_26;
begin
n1 <= s29_1(9 downto 9);
n2 <= s25_1 & s25_2;
process (clock_c) begin
  if rising_edge(clock_c) then
    if i5 = "1" then
      n3 <= "0";
    elsif i4 = "1" then
      n3 <= s29_2;
    end if;
  end if;
end process;
process (clock_c) begin
  if rising_edge(clock_c) then
    if i5 = "1" then
      n4 <= "0";
    elsif i4 = "1" then
      n4 <= n3;
    end if;
  end if;
end process;
process (clock_c) begin
  if rising_edge(clock_c) then
    if i5 = "1" then
      n5 <= "0";
    elsif i4 = "1" then
      n5 <= n4;
    end if;
  end if;
end process;
process (clock_c) begin
  if rising_edge(clock_c) then
    if i5 = "1" then
      n6 <= "0";
    elsif i4 = "1" then
      n6 <= n5;
    end if;
  end if;
end process;
n7 <= s29_1(9 downto 9) &
  s29_1(8 downto 8) &
  s29_1(7 downto 7) &
  s29_1(6 downto 6) &
  s29_1(5 downto 5) &
  s29_1(4 downto 4) &
  s29_1(3 downto 3) &
  s29_1(2 downto 2) &
  s29_1(1 downto 1);
process (clock_c) begin
  if rising_edge(clock_c) then
    if i5 = "1" then
      n8 <= "000000000";
    elsif i4 = "1" then
      n8 <= n7;
    end if;
  end if;
end process;
process (clock_c) begin
  if rising_edge(clock_c) then
    if i5 = "1" then
      n9 <= "000000000";
    elsif i4 = "1" then
      n9 <= n8;
    end if;
  end if;
end process;
process (clock_c) begin
  if rising_edge(clock_c) then
    if i5 = "1" then
      n10 <= "000000000";
    elsif i4 = "1" then
      n10 <= n9;
    end if;
  end if;
end process;
process (clock_c) begin
  if rising_edge(clock_c) then
    if i5 = "1" then
      n11 <= "000000000";
    elsif i4 = "1" then
      n11 <= n10;
    end if;
  end if;
end process;
n12 <= s29_1(0 downto 0);
process (clock_c) begin
  if rising_edge(clock_c) then
    if i5 = "1" then
      n13 <= "0";
    elsif i4 = "1" then
      n13 <= n12;
    end if;
  end if;
end process;
process (clock_c) begin
  if rising_edge(clock_c) then
    if i5 = "1" then
      n14 <= "0";
    elsif i4 = "1" then
      n14 <= n13;
    end if;
  end if;
end process;
process (clock_c) begin
  if rising_edge(clock_c) then
    if i5 = "1" then
      n15 <= "0";
    elsif i4 = "1" then
      n15 <= n14;
    end if;
  end if;
end process;
process (clock_c) begin
  if rising_edge(clock_c) then
    if i5 = "1" then
      n16 <= "0";
    elsif i4 = "1" then
      n16 <= n15;
    end if;
  end if;
end process;
n17 <= not n16;
n18 <= s28_2 & s28_1;
n19 <= s28_3(63 downto 63) &
  s28_3(62 downto 62) &
  s28_3(61 downto 61) &
  s28_3(60 downto 60) &
  s28_3(59 downto 59) &
  s28_3(58 downto 58) &
  s28_3(57 downto 57) &
  s28_3(56 downto 56) &
  s28_3(55 downto 55) &
  s28_3(54 downto 54) &
  s28_3(53 downto 53) &
  s28_3(52 downto 52) &
  s28_3(51 downto 51) &
  s28_3(50 downto 50) &
  s28_3(49 downto 49) &
  s28_3(48 downto 48) &
  s28_3(47 downto 47) &
  s28_3(46 downto 46) &
  s28_3(45 downto 45) &
  s28_3(44 downto 44) &
  s28_3(43 downto 43) &
  s28_3(42 downto 42) &
  s28_3(41 downto 41) &
  s28_3(40 downto 40) &
  s28_3(39 downto 39) &
  s28_3(38 downto 38) &
  s28_3(37 downto 37) &
  s28_3(36 downto 36) &
  s28_3(35 downto 35) &
  s28_3(34 downto 34) &
  s28_3(33 downto 33) &
  s28_3(32 downto 32);
n20 <= s28_3(31 downto 31) &
  s28_3(30 downto 30) &
  s28_3(29 downto 29) &
  s28_3(28 downto 28) &
  s28_3(27 downto 27) &
  s28_3(26 downto 26) &
  s28_3(25 downto 25) &
  s28_3(24 downto 24) &
  s28_3(23 downto 23) &
  s28_3(22 downto 22) &
  s28_3(21 downto 21) &
  s28_3(20 downto 20) &
  s28_3(19 downto 19) &
  s28_3(18 downto 18) &
  s28_3(17 downto 17) &
  s28_3(16 downto 16) &
  s28_3(15 downto 15) &
  s28_3(14 downto 14) &
  s28_3(13 downto 13) &
  s28_3(12 downto 12) &
  s28_3(11 downto 11) &
  s28_3(10 downto 10) &
  s28_3(9 downto 9) &
  s28_3(8 downto 8) &
  s28_3(7 downto 7) &
  s28_3(6 downto 6) &
  s28_3(5 downto 5) &
  s28_3(4 downto 4) &
  s28_3(3 downto 3) &
  s28_3(2 downto 2) &
  s28_3(1 downto 1) &
  s28_3(0 downto 0);
n21 <= s27_1(63 downto 63) &
  s27_1(62 downto 62) &
  s27_1(61 downto 61) &
  s27_1(60 downto 60) &
  s27_1(59 downto 59) &
  s27_1(58 downto 58) &
  s27_1(57 downto 57) &
  s27_1(56 downto 56) &
  s27_1(55 downto 55) &
  s27_1(54 downto 54) &
  s27_1(53 downto 53) &
  s27_1(52 downto 52) &
  s27_1(51 downto 51) &
  s27_1(50 downto 50) &
  s27_1(49 downto 49) &
  s27_1(48 downto 48) &
  s27_1(47 downto 47) &
  s27_1(46 downto 46) &
  s27_1(45 downto 45) &
  s27_1(44 downto 44) &
  s27_1(43 downto 43) &
  s27_1(42 downto 42) &
  s27_1(41 downto 41) &
  s27_1(40 downto 40) &
  s27_1(39 downto 39) &
  s27_1(38 downto 38) &
  s27_1(37 downto 37) &
  s27_1(36 downto 36) &
  s27_1(35 downto 35) &
  s27_1(34 downto 34) &
  s27_1(33 downto 33) &
  s27_1(32 downto 32);
n22 <= s27_1(31 downto 31) &
  s27_1(30 downto 30) &
  s27_1(29 downto 29) &
  s27_1(28 downto 28) &
  s27_1(27 downto 27) &
  s27_1(26 downto 26) &
  s27_1(25 downto 25) &
  s27_1(24 downto 24) &
  s27_1(23 downto 23) &
  s27_1(22 downto 22) &
  s27_1(21 downto 21) &
  s27_1(20 downto 20) &
  s27_1(19 downto 19) &
  s27_1(18 downto 18) &
  s27_1(17 downto 17) &
  s27_1(16 downto 16) &
  s27_1(15 downto 15) &
  s27_1(14 downto 14) &
  s27_1(13 downto 13) &
  s27_1(12 downto 12) &
  s27_1(11 downto 11) &
  s27_1(10 downto 10) &
  s27_1(9 downto 9) &
  s27_1(8 downto 8) &
  s27_1(7 downto 7) &
  s27_1(6 downto 6) &
  s27_1(5 downto 5) &
  s27_1(4 downto 4) &
  s27_1(3 downto 3) &
  s27_1(2 downto 2) &
  s27_1(1 downto 1) &
  s27_1(0 downto 0);
n23 <= n20 when s26_1 = "1" else n19;
n24 <= n22 when s26_1 = "1" else n21;
s25 : cf_fft_2048_16_7 port map (clock_c, i2, i3, n1, i4, i5, s25_1, s25_2);
s26 : cf_fft_2048_16_35 port map (clock_c, n18, i4, i5, s26_1);
s27 : cf_fft_2048_16_31 port map (clock_c, n2, n6, n11, n16, i4, i5, s27_1);
s28 : cf_fft_2048_16_30 port map (clock_c, n2, n6, n11, n17, i4, i5, s28_1, s28_2, s28_3);
s29 : cf_fft_2048_16_26 port map (clock_c, i1, i4, i5, s29_1, s29_2);
o3 <= n24;
o2 <= n23;
o1 <= s28_1;
end architecture rtl;

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
entity cf_fft_2048_16_5 is
port (
clock_c : in std_logic;
i1 : in  unsigned(0 downto 0);
i2 : in  unsigned(31 downto 0);
i3 : in  unsigned(31 downto 0);
i4 : in  unsigned(0 downto 0);
i5 : in  unsigned(0 downto 0);
o1 : out unsigned(0 downto 0);
o2 : out unsigned(31 downto 0);
o3 : out unsigned(31 downto 0));
end entity cf_fft_2048_16_5;
architecture rtl of cf_fft_2048_16_5 is
signal n1 : unsigned(0 downto 0);
signal n2 : unsigned(63 downto 0);
signal n3 : unsigned(0 downto 0) := "0";
signal n4 : unsigned(0 downto 0) := "0";
signal n5 : unsigned(0 downto 0) := "0";
signal n6 : unsigned(0 downto 0) := "0";
signal n7 : unsigned(8 downto 0);
signal n8 : unsigned(8 downto 0) := "000000000";
signal n9 : unsigned(8 downto 0) := "000000000";
signal n10 : unsigned(8 downto 0) := "000000000";
signal n11 : unsigned(8 downto 0) := "000000000";
signal n12 : unsigned(0 downto 0);
signal n13 : unsigned(0 downto 0) := "0";
signal n14 : unsigned(0 downto 0) := "0";
signal n15 : unsigned(0 downto 0) := "0";
signal n16 : unsigned(0 downto 0) := "0";
signal n17 : unsigned(0 downto 0);
signal n18 : unsigned(1 downto 0);
signal n19 : unsigned(31 downto 0);
signal n20 : unsigned(31 downto 0);
signal n21 : unsigned(31 downto 0);
signal n22 : unsigned(31 downto 0);
signal n23 : unsigned(31 downto 0);
signal n24 : unsigned(31 downto 0);
signal s25_1 : unsigned(31 downto 0);
signal s25_2 : unsigned(31 downto 0);
signal s26_1 : unsigned(0 downto 0);
signal s27_1 : unsigned(63 downto 0);
signal s28_1 : unsigned(0 downto 0);
signal s28_2 : unsigned(0 downto 0);
signal s28_3 : unsigned(63 downto 0);
signal s29_1 : unsigned(9 downto 0);
signal s29_2 : unsigned(0 downto 0);
component cf_fft_2048_16_7 is
port (
clock_c : in std_logic;
i1 : in  unsigned(31 downto 0);
i2 : in  unsigned(31 downto 0);
i3 : in  unsigned(0 downto 0);
i4 : in  unsigned(0 downto 0);
i5 : in  unsigned(0 downto 0);
o1 : out unsigned(31 downto 0);
o2 : out unsigned(31 downto 0));
end component cf_fft_2048_16_7;
component cf_fft_2048_16_35 is
port (
clock_c : in std_logic;
i1 : in  unsigned(1 downto 0);
i2 : in  unsigned(0 downto 0);
i3 : in  unsigned(0 downto 0);
o1 : out unsigned(0 downto 0));
end component cf_fft_2048_16_35;
component cf_fft_2048_16_31 is
port (
clock_c : in std_logic;
i1 : in  unsigned(63 downto 0);
i2 : in  unsigned(0 downto 0);
i3 : in  unsigned(8 downto 0);
i4 : in  unsigned(0 downto 0);
i5 : in  unsigned(0 downto 0);
i6 : in  unsigned(0 downto 0);
o1 : out unsigned(63 downto 0));
end component cf_fft_2048_16_31;
component cf_fft_2048_16_30 is
port (
clock_c : in std_logic;
i1 : in  unsigned(63 downto 0);
i2 : in  unsigned(0 downto 0);
i3 : in  unsigned(8 downto 0);
i4 : in  unsigned(0 downto 0);
i5 : in  unsigned(0 downto 0);
i6 : in  unsigned(0 downto 0);
o1 : out unsigned(0 downto 0);
o2 : out unsigned(0 downto 0);
o3 : out unsigned(63 downto 0));
end component cf_fft_2048_16_30;
component cf_fft_2048_16_26 is
port (
clock_c : in std_logic;
i1 : in  unsigned(0 downto 0);
i2 : in  unsigned(0 downto 0);
i3 : in  unsigned(0 downto 0);
o1 : out unsigned(9 downto 0);
o2 : out unsigned(0 downto 0));
end component cf_fft_2048_16_26;
begin
n1 <= "0";
n2 <= s25_1 & s25_2;
process (clock_c) begin
  if rising_edge(clock_c) then
    if i5 = "1" then
      n3 <= "0";
    elsif i4 = "1" then
      n3 <= s29_2;
    end if;
  end if;
end process;
process (clock_c) begin
  if rising_edge(clock_c) then
    if i5 = "1" then
      n4 <= "0";
    elsif i4 = "1" then
      n4 <= n3;
    end if;
  end if;
end process;
process (clock_c) begin
  if rising_edge(clock_c) then
    if i5 = "1" then
      n5 <= "0";
    elsif i4 = "1" then
      n5 <= n4;
    end if;
  end if;
end process;
process (clock_c) begin
  if rising_edge(clock_c) then
    if i5 = "1" then
      n6 <= "0";
    elsif i4 = "1" then
      n6 <= n5;
    end if;
  end if;
end process;
n7 <= s29_1(9 downto 9) &
  s29_1(8 downto 8) &
  s29_1(7 downto 7) &
  s29_1(6 downto 6) &
  s29_1(5 downto 5) &
  s29_1(4 downto 4) &
  s29_1(3 downto 3) &
  s29_1(2 downto 2) &
  s29_1(1 downto 1);
process (clock_c) begin
  if rising_edge(clock_c) then
    if i5 = "1" then
      n8 <= "000000000";
    elsif i4 = "1" then
      n8 <= n7;
    end if;
  end if;
end process;
process (clock_c) begin
  if rising_edge(clock_c) then
    if i5 = "1" then
      n9 <= "000000000";
    elsif i4 = "1" then
      n9 <= n8;
    end if;
  end if;
end process;
process (clock_c) begin
  if rising_edge(clock_c) then
    if i5 = "1" then
      n10 <= "000000000";
    elsif i4 = "1" then
      n10 <= n9;
    end if;
  end if;
end process;
process (clock_c) begin
  if rising_edge(clock_c) then
    if i5 = "1" then
      n11 <= "000000000";
    elsif i4 = "1" then
      n11 <= n10;
    end if;
  end if;
end process;
n12 <= s29_1(0 downto 0);
process (clock_c) begin
  if rising_edge(clock_c) then
    if i5 = "1" then
      n13 <= "0";
    elsif i4 = "1" then
      n13 <= n12;
    end if;
  end if;
end process;
process (clock_c) begin
  if rising_edge(clock_c) then
    if i5 = "1" then
      n14 <= "0";
    elsif i4 = "1" then
      n14 <= n13;
    end if;
  end if;
end process;
process (clock_c) begin
  if rising_edge(clock_c) then
    if i5 = "1" then
      n15 <= "0";
    elsif i4 = "1" then
      n15 <= n14;
    end if;
  end if;
end process;
process (clock_c) begin
  if rising_edge(clock_c) then
    if i5 = "1" then
      n16 <= "0";
    elsif i4 = "1" then
      n16 <= n15;
    end if;
  end if;
end process;
n17 <= not n16;
n18 <= s28_2 & s28_1;
n19 <= s28_3(63 downto 63) &
  s28_3(62 downto 62) &
  s28_3(61 downto 61) &
  s28_3(60 downto 60) &
  s28_3(59 downto 59) &
  s28_3(58 downto 58) &
  s28_3(57 downto 57) &
  s28_3(56 downto 56) &
  s28_3(55 downto 55) &
  s28_3(54 downto 54) &
  s28_3(53 downto 53) &
  s28_3(52 downto 52) &
  s28_3(51 downto 51) &
  s28_3(50 downto 50) &
  s28_3(49 downto 49) &
  s28_3(48 downto 48) &
  s28_3(47 downto 47) &
  s28_3(46 downto 46) &
  s28_3(45 downto 45) &
  s28_3(44 downto 44) &
  s28_3(43 downto 43) &
  s28_3(42 downto 42) &
  s28_3(41 downto 41) &
  s28_3(40 downto 40) &
  s28_3(39 downto 39) &
  s28_3(38 downto 38) &
  s28_3(37 downto 37) &
  s28_3(36 downto 36) &
  s28_3(35 downto 35) &
  s28_3(34 downto 34) &
  s28_3(33 downto 33) &
  s28_3(32 downto 32);
n20 <= s28_3(31 downto 31) &
  s28_3(30 downto 30) &
  s28_3(29 downto 29) &
  s28_3(28 downto 28) &
  s28_3(27 downto 27) &
  s28_3(26 downto 26) &
  s28_3(25 downto 25) &
  s28_3(24 downto 24) &
  s28_3(23 downto 23) &
  s28_3(22 downto 22) &
  s28_3(21 downto 21) &
  s28_3(20 downto 20) &
  s28_3(19 downto 19) &
  s28_3(18 downto 18) &
  s28_3(17 downto 17) &
  s28_3(16 downto 16) &
  s28_3(15 downto 15) &
  s28_3(14 downto 14) &
  s28_3(13 downto 13) &
  s28_3(12 downto 12) &
  s28_3(11 downto 11) &
  s28_3(10 downto 10) &
  s28_3(9 downto 9) &
  s28_3(8 downto 8) &
  s28_3(7 downto 7) &
  s28_3(6 downto 6) &
  s28_3(5 downto 5) &
  s28_3(4 downto 4) &
  s28_3(3 downto 3) &
  s28_3(2 downto 2) &
  s28_3(1 downto 1) &
  s28_3(0 downto 0);
n21 <= s27_1(63 downto 63) &
  s27_1(62 downto 62) &
  s27_1(61 downto 61) &
  s27_1(60 downto 60) &
  s27_1(59 downto 59) &
  s27_1(58 downto 58) &
  s27_1(57 downto 57) &
  s27_1(56 downto 56) &
  s27_1(55 downto 55) &
  s27_1(54 downto 54) &
  s27_1(53 downto 53) &
  s27_1(52 downto 52) &
  s27_1(51 downto 51) &
  s27_1(50 downto 50) &
  s27_1(49 downto 49) &
  s27_1(48 downto 48) &
  s27_1(47 downto 47) &
  s27_1(46 downto 46) &
  s27_1(45 downto 45) &
  s27_1(44 downto 44) &
  s27_1(43 downto 43) &
  s27_1(42 downto 42) &
  s27_1(41 downto 41) &
  s27_1(40 downto 40) &
  s27_1(39 downto 39) &
  s27_1(38 downto 38) &
  s27_1(37 downto 37) &
  s27_1(36 downto 36) &
  s27_1(35 downto 35) &
  s27_1(34 downto 34) &
  s27_1(33 downto 33) &
  s27_1(32 downto 32);
n22 <= s27_1(31 downto 31) &
  s27_1(30 downto 30) &
  s27_1(29 downto 29) &
  s27_1(28 downto 28) &
  s27_1(27 downto 27) &
  s27_1(26 downto 26) &
  s27_1(25 downto 25) &
  s27_1(24 downto 24) &
  s27_1(23 downto 23) &
  s27_1(22 downto 22) &
  s27_1(21 downto 21) &
  s27_1(20 downto 20) &
  s27_1(19 downto 19) &
  s27_1(18 downto 18) &
  s27_1(17 downto 17) &
  s27_1(16 downto 16) &
  s27_1(15 downto 15) &
  s27_1(14 downto 14) &
  s27_1(13 downto 13) &
  s27_1(12 downto 12) &
  s27_1(11 downto 11) &
  s27_1(10 downto 10) &
  s27_1(9 downto 9) &
  s27_1(8 downto 8) &
  s27_1(7 downto 7) &
  s27_1(6 downto 6) &
  s27_1(5 downto 5) &
  s27_1(4 downto 4) &
  s27_1(3 downto 3) &
  s27_1(2 downto 2) &
  s27_1(1 downto 1) &
  s27_1(0 downto 0);
n23 <= n20 when s26_1 = "1" else n19;
n24 <= n22 when s26_1 = "1" else n21;
s25 : cf_fft_2048_16_7 port map (clock_c, i2, i3, n1, i4, i5, s25_1, s25_2);
s26 : cf_fft_2048_16_35 port map (clock_c, n18, i4, i5, s26_1);
s27 : cf_fft_2048_16_31 port map (clock_c, n2, n6, n11, n16, i4, i5, s27_1);
s28 : cf_fft_2048_16_30 port map (clock_c, n2, n6, n11, n17, i4, i5, s28_1, s28_2, s28_3);
s29 : cf_fft_2048_16_26 port map (clock_c, i1, i4, i5, s29_1, s29_2);
o3 <= n24;
o2 <= n23;
o1 <= s28_1;
end architecture rtl;

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
entity cf_fft_2048_16_4 is
port (
clock_c : in std_logic;
i1 : in  unsigned(0 downto 0);
i2 : in  unsigned(63 downto 0);
i3 : in  unsigned(0 downto 0);
i4 : in  unsigned(8 downto 0);
i5 : in  unsigned(0 downto 0);
i6 : in  unsigned(0 downto 0);
o1 : out unsigned(63 downto 0));
end entity cf_fft_2048_16_4;
architecture rtl of cf_fft_2048_16_4 is
signal n1 : unsigned(8 downto 0);
signal n2 : unsigned(8 downto 0);
signal n3 : unsigned(8 downto 0) := "000000000";
signal n4 : unsigned(0 downto 0);
signal n5 : unsigned(0 downto 0);
signal n6 : unsigned(63 downto 0);
signal n6a : unsigned(8 downto 0) := "000000000";
type   n6mt is array (511 downto 0) of unsigned(63 downto 0);
signal n6m : n6mt;
signal n7 : unsigned(0 downto 0);
signal n8 : unsigned(63 downto 0);
signal n8a : unsigned(8 downto 0) := "000000000";
type   n8mt is array (511 downto 0) of unsigned(63 downto 0);
signal n8m : n8mt;
signal n9 : unsigned(0 downto 0) := "0";
signal n10 : unsigned(63 downto 0);
signal n11 : unsigned(0 downto 0);
signal s12_1 : unsigned(0 downto 0);
component cf_fft_2048_16_32 is
port (
clock_c : in std_logic;
i1 : in  unsigned(0 downto 0);
i2 : in  unsigned(0 downto 0);
i3 : in  unsigned(0 downto 0);
o1 : out unsigned(0 downto 0));
end component cf_fft_2048_16_32;
begin
n1 <= "000000001";
n2 <= n3 + n1;
process (clock_c) begin
  if rising_edge(clock_c) then
    if n11 = "1" then
      n3 <= "000000000";
    elsif i5 = "1" then
      n3 <= n2;
    end if;
  end if;
end process;
n4 <= not s12_1;
n5 <= i3 and n4;
process (clock_c) begin
  if rising_edge(clock_c) then
    if i5 = "1" then
      if n5 = "1" then
        n6m(to_integer(i4)) <= i2;
      end if;
      n6a <= n3;
    end if;
  end if;
end process;
n6 <= n6m(to_integer(n6a));
n7 <= i3 and s12_1;
process (clock_c) begin
  if rising_edge(clock_c) then
    if i5 = "1" then
      if n7 = "1" then
        n8m(to_integer(i4)) <= i2;
      end if;
      n8a <= n3;
    end if;
  end if;
end process;
n8 <= n8m(to_integer(n8a));
process (clock_c) begin
  if rising_edge(clock_c) then
    if i6 = "1" then
      n9 <= "0";
    elsif i5 = "1" then
      n9 <= n4;
    end if;
  end if;
end process;
n10 <= n8 when n9 = "1" else n6;
n11 <= i1 or i6;
s12 : cf_fft_2048_16_32 port map (clock_c, i1, i5, i6, s12_1);
o1 <= n10;
end architecture rtl;

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
entity cf_fft_2048_16_3 is
port (
clock_c : in std_logic;
i1 : in  unsigned(0 downto 0);
i2 : in  unsigned(63 downto 0);
i3 : in  unsigned(0 downto 0);
i4 : in  unsigned(8 downto 0);
i5 : in  unsigned(0 downto 0);
i6 : in  unsigned(0 downto 0);
o1 : out unsigned(0 downto 0);
o2 : out unsigned(0 downto 0);
o3 : out unsigned(63 downto 0));
end entity cf_fft_2048_16_3;
architecture rtl of cf_fft_2048_16_3 is
signal n1 : unsigned(8 downto 0);
signal n2 : unsigned(8 downto 0);
signal n3 : unsigned(8 downto 0) := "000000000";
signal n4 : unsigned(0 downto 0);
signal n5 : unsigned(0 downto 0) := "0";
signal n6 : unsigned(8 downto 0);
signal n7 : unsigned(0 downto 0);
signal n8 : unsigned(0 downto 0);
signal n9 : unsigned(63 downto 0);
signal n9a : unsigned(8 downto 0) := "000000000";
type   n9mt is array (511 downto 0) of unsigned(63 downto 0);
signal n9m : n9mt;
signal n10 : unsigned(0 downto 0);
signal n11 : unsigned(63 downto 0);
signal n11a : unsigned(8 downto 0) := "000000000";
type   n11mt is array (511 downto 0) of unsigned(63 downto 0);
signal n11m : n11mt;
signal n12 : unsigned(0 downto 0) := "0";
signal n13 : unsigned(63 downto 0);
signal n14 : unsigned(0 downto 0);
signal s15_1 : unsigned(0 downto 0);
component cf_fft_2048_16_32 is
port (
clock_c : in std_logic;
i1 : in  unsigned(0 downto 0);
i2 : in  unsigned(0 downto 0);
i3 : in  unsigned(0 downto 0);
o1 : out unsigned(0 downto 0));
end component cf_fft_2048_16_32;
begin
n1 <= "000000001";
n2 <= n3 + n1;
process (clock_c) begin
  if rising_edge(clock_c) then
    if n14 = "1" then
      n3 <= "000000000";
    elsif i5 = "1" then
      n3 <= n2;
    end if;
  end if;
end process;
n4 <= not s15_1;
process (clock_c) begin
  if rising_edge(clock_c) then
    if i6 = "1" then
      n5 <= "0";
    elsif i5 = "1" then
      n5 <= i1;
    end if;
  end if;
end process;
n6 <= "000000000";
n7 <= "1" when n3 = n6 else "0";
n8 <= i3 and n4;
process (clock_c) begin
  if rising_edge(clock_c) then
    if i5 = "1" then
      if n8 = "1" then
        n9m(to_integer(i4)) <= i2;
      end if;
      n9a <= n3;
    end if;
  end if;
end process;
n9 <= n9m(to_integer(n9a));
n10 <= i3 and s15_1;
process (clock_c) begin
  if rising_edge(clock_c) then
    if i5 = "1" then
      if n10 = "1" then
        n11m(to_integer(i4)) <= i2;
      end if;
      n11a <= n3;
    end if;
  end if;
end process;
n11 <= n11m(to_integer(n11a));
process (clock_c) begin
  if rising_edge(clock_c) then
    if i6 = "1" then
      n12 <= "0";
    elsif i5 = "1" then
      n12 <= n4;
    end if;
  end if;
end process;
n13 <= n11 when n12 = "1" else n9;
n14 <= i1 or i6;
s15 : cf_fft_2048_16_32 port map (clock_c, i1, i5, i6, s15_1);
o3 <= n13;
o2 <= n7;
o1 <= n5;
end architecture rtl;

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
entity cf_fft_2048_16_2 is
port (
clock_c : in std_logic;
i1 : in  unsigned(0 downto 0);
i2 : in  unsigned(31 downto 0);
i3 : in  unsigned(31 downto 0);
i4 : in  unsigned(0 downto 0);
i5 : in  unsigned(0 downto 0);
o1 : out unsigned(0 downto 0);
o2 : out unsigned(31 downto 0);
o3 : out unsigned(31 downto 0));
end entity cf_fft_2048_16_2;
architecture rtl of cf_fft_2048_16_2 is
signal n1 : unsigned(63 downto 0);
signal n2 : unsigned(0 downto 0);
signal n3 : unsigned(0 downto 0);
signal n4 : unsigned(8 downto 0);
signal n5 : unsigned(8 downto 0);
signal n6 : unsigned(1 downto 0);
signal n7 : unsigned(31 downto 0);
signal n8 : unsigned(31 downto 0);
signal n9 : unsigned(31 downto 0);
signal n10 : unsigned(31 downto 0);
signal n11 : unsigned(31 downto 0);
signal n12 : unsigned(31 downto 0);
signal s13_1 : unsigned(0 downto 0);
signal s14_1 : unsigned(63 downto 0);
signal s15_1 : unsigned(0 downto 0);
signal s15_2 : unsigned(0 downto 0);
signal s15_3 : unsigned(63 downto 0);
signal s16_1 : unsigned(9 downto 0);
signal s16_2 : unsigned(0 downto 0);
component cf_fft_2048_16_35 is
port (
clock_c : in std_logic;
i1 : in  unsigned(1 downto 0);
i2 : in  unsigned(0 downto 0);
i3 : in  unsigned(0 downto 0);
o1 : out unsigned(0 downto 0));
end component cf_fft_2048_16_35;
component cf_fft_2048_16_4 is
port (
clock_c : in std_logic;
i1 : in  unsigned(0 downto 0);
i2 : in  unsigned(63 downto 0);
i3 : in  unsigned(0 downto 0);
i4 : in  unsigned(8 downto 0);
i5 : in  unsigned(0 downto 0);
i6 : in  unsigned(0 downto 0);
o1 : out unsigned(63 downto 0));
end component cf_fft_2048_16_4;
component cf_fft_2048_16_3 is
port (
clock_c : in std_logic;
i1 : in  unsigned(0 downto 0);
i2 : in  unsigned(63 downto 0);
i3 : in  unsigned(0 downto 0);
i4 : in  unsigned(8 downto 0);
i5 : in  unsigned(0 downto 0);
i6 : in  unsigned(0 downto 0);
o1 : out unsigned(0 downto 0);
o2 : out unsigned(0 downto 0);
o3 : out unsigned(63 downto 0));
end component cf_fft_2048_16_3;
component cf_fft_2048_16_26 is
port (
clock_c : in std_logic;
i1 : in  unsigned(0 downto 0);
i2 : in  unsigned(0 downto 0);
i3 : in  unsigned(0 downto 0);
o1 : out unsigned(9 downto 0);
o2 : out unsigned(0 downto 0));
end component cf_fft_2048_16_26;
begin
n1 <= i2 & i3;
n2 <= s16_1(9 downto 9);
n3 <= not n2;
n4 <= s16_1(8 downto 8) &
  s16_1(7 downto 7) &
  s16_1(6 downto 6) &
  s16_1(5 downto 5) &
  s16_1(4 downto 4) &
  s16_1(3 downto 3) &
  s16_1(2 downto 2) &
  s16_1(1 downto 1) &
  s16_1(0 downto 0);
n5 <= n4(0 downto 0) &
  n4(1 downto 1) &
  n4(2 downto 2) &
  n4(3 downto 3) &
  n4(4 downto 4) &
  n4(5 downto 5) &
  n4(6 downto 6) &
  n4(7 downto 7) &
  n4(8 downto 8);
n6 <= s15_2 & s15_1;
n7 <= s15_3(63 downto 63) &
  s15_3(62 downto 62) &
  s15_3(61 downto 61) &
  s15_3(60 downto 60) &
  s15_3(59 downto 59) &
  s15_3(58 downto 58) &
  s15_3(57 downto 57) &
  s15_3(56 downto 56) &
  s15_3(55 downto 55) &
  s15_3(54 downto 54) &
  s15_3(53 downto 53) &
  s15_3(52 downto 52) &
  s15_3(51 downto 51) &
  s15_3(50 downto 50) &
  s15_3(49 downto 49) &
  s15_3(48 downto 48) &
  s15_3(47 downto 47) &
  s15_3(46 downto 46) &
  s15_3(45 downto 45) &
  s15_3(44 downto 44) &
  s15_3(43 downto 43) &
  s15_3(42 downto 42) &
  s15_3(41 downto 41) &
  s15_3(40 downto 40) &
  s15_3(39 downto 39) &
  s15_3(38 downto 38) &
  s15_3(37 downto 37) &
  s15_3(36 downto 36) &
  s15_3(35 downto 35) &
  s15_3(34 downto 34) &
  s15_3(33 downto 33) &
  s15_3(32 downto 32);
n8 <= s15_3(31 downto 31) &
  s15_3(30 downto 30) &
  s15_3(29 downto 29) &
  s15_3(28 downto 28) &
  s15_3(27 downto 27) &
  s15_3(26 downto 26) &
  s15_3(25 downto 25) &
  s15_3(24 downto 24) &
  s15_3(23 downto 23) &
  s15_3(22 downto 22) &
  s15_3(21 downto 21) &
  s15_3(20 downto 20) &
  s15_3(19 downto 19) &
  s15_3(18 downto 18) &
  s15_3(17 downto 17) &
  s15_3(16 downto 16) &
  s15_3(15 downto 15) &
  s15_3(14 downto 14) &
  s15_3(13 downto 13) &
  s15_3(12 downto 12) &
  s15_3(11 downto 11) &
  s15_3(10 downto 10) &
  s15_3(9 downto 9) &
  s15_3(8 downto 8) &
  s15_3(7 downto 7) &
  s15_3(6 downto 6) &
  s15_3(5 downto 5) &
  s15_3(4 downto 4) &
  s15_3(3 downto 3) &
  s15_3(2 downto 2) &
  s15_3(1 downto 1) &
  s15_3(0 downto 0);
n9 <= s14_1(63 downto 63) &
  s14_1(62 downto 62) &
  s14_1(61 downto 61) &
  s14_1(60 downto 60) &
  s14_1(59 downto 59) &
  s14_1(58 downto 58) &
  s14_1(57 downto 57) &
  s14_1(56 downto 56) &
  s14_1(55 downto 55) &
  s14_1(54 downto 54) &
  s14_1(53 downto 53) &
  s14_1(52 downto 52) &
  s14_1(51 downto 51) &
  s14_1(50 downto 50) &
  s14_1(49 downto 49) &
  s14_1(48 downto 48) &
  s14_1(47 downto 47) &
  s14_1(46 downto 46) &
  s14_1(45 downto 45) &
  s14_1(44 downto 44) &
  s14_1(43 downto 43) &
  s14_1(42 downto 42) &
  s14_1(41 downto 41) &
  s14_1(40 downto 40) &
  s14_1(39 downto 39) &
  s14_1(38 downto 38) &
  s14_1(37 downto 37) &
  s14_1(36 downto 36) &
  s14_1(35 downto 35) &
  s14_1(34 downto 34) &
  s14_1(33 downto 33) &
  s14_1(32 downto 32);
n10 <= s14_1(31 downto 31) &
  s14_1(30 downto 30) &
  s14_1(29 downto 29) &
  s14_1(28 downto 28) &
  s14_1(27 downto 27) &
  s14_1(26 downto 26) &
  s14_1(25 downto 25) &
  s14_1(24 downto 24) &
  s14_1(23 downto 23) &
  s14_1(22 downto 22) &
  s14_1(21 downto 21) &
  s14_1(20 downto 20) &
  s14_1(19 downto 19) &
  s14_1(18 downto 18) &
  s14_1(17 downto 17) &
  s14_1(16 downto 16) &
  s14_1(15 downto 15) &
  s14_1(14 downto 14) &
  s14_1(13 downto 13) &
  s14_1(12 downto 12) &
  s14_1(11 downto 11) &
  s14_1(10 downto 10) &
  s14_1(9 downto 9) &
  s14_1(8 downto 8) &
  s14_1(7 downto 7) &
  s14_1(6 downto 6) &
  s14_1(5 downto 5) &
  s14_1(4 downto 4) &
  s14_1(3 downto 3) &
  s14_1(2 downto 2) &
  s14_1(1 downto 1) &
  s14_1(0 downto 0);
n11 <= n8 when s13_1 = "1" else n7;
n12 <= n10 when s13_1 = "1" else n9;
s13 : cf_fft_2048_16_35 port map (clock_c, n6, i4, i5, s13_1);
s14 : cf_fft_2048_16_4 port map (clock_c, s16_2, n1, n2, n5, i4, i5, s14_1);
s15 : cf_fft_2048_16_3 port map (clock_c, s16_2, n1, n3, n5, i4, i5, s15_1, s15_2, s15_3);
s16 : cf_fft_2048_16_26 port map (clock_c, i1, i4, i5, s16_1, s16_2);
o3 <= n12;
o2 <= n11;
o1 <= s15_1;
end architecture rtl;

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
entity cf_fft_2048_16_1 is
port (
clock_c : in std_logic;
i1 : in  unsigned(0 downto 0);
i2 : in  unsigned(31 downto 0);
i3 : in  unsigned(31 downto 0);
i4 : in  unsigned(0 downto 0);
i5 : in  unsigned(0 downto 0);
o1 : out unsigned(0 downto 0);
o2 : out unsigned(31 downto 0);
o3 : out unsigned(31 downto 0));
end entity cf_fft_2048_16_1;
architecture rtl of cf_fft_2048_16_1 is
signal s1_1 : unsigned(0 downto 0);
signal s1_2 : unsigned(31 downto 0);
signal s1_3 : unsigned(31 downto 0);
signal s2_1 : unsigned(0 downto 0);
signal s2_2 : unsigned(31 downto 0);
signal s2_3 : unsigned(31 downto 0);
signal s3_1 : unsigned(0 downto 0);
signal s3_2 : unsigned(31 downto 0);
signal s3_3 : unsigned(31 downto 0);
signal s4_1 : unsigned(0 downto 0);
signal s4_2 : unsigned(31 downto 0);
signal s4_3 : unsigned(31 downto 0);
signal s5_1 : unsigned(0 downto 0);
signal s5_2 : unsigned(31 downto 0);
signal s5_3 : unsigned(31 downto 0);
component cf_fft_2048_16_25 is
port (
clock_c : in std_logic;
i1 : in  unsigned(0 downto 0);
i2 : in  unsigned(31 downto 0);
i3 : in  unsigned(31 downto 0);
i4 : in  unsigned(0 downto 0);
i5 : in  unsigned(0 downto 0);
o1 : out unsigned(0 downto 0);
o2 : out unsigned(31 downto 0);
o3 : out unsigned(31 downto 0));
end component cf_fft_2048_16_25;
component cf_fft_2048_16_8 is
port (
clock_c : in std_logic;
i1 : in  unsigned(0 downto 0);
i2 : in  unsigned(31 downto 0);
i3 : in  unsigned(31 downto 0);
i4 : in  unsigned(0 downto 0);
i5 : in  unsigned(0 downto 0);
o1 : out unsigned(0 downto 0);
o2 : out unsigned(31 downto 0);
o3 : out unsigned(31 downto 0));
end component cf_fft_2048_16_8;
component cf_fft_2048_16_6 is
port (
clock_c : in std_logic;
i1 : in  unsigned(0 downto 0);
i2 : in  unsigned(31 downto 0);
i3 : in  unsigned(31 downto 0);
i4 : in  unsigned(0 downto 0);
i5 : in  unsigned(0 downto 0);
o1 : out unsigned(0 downto 0);
o2 : out unsigned(31 downto 0);
o3 : out unsigned(31 downto 0));
end component cf_fft_2048_16_6;
component cf_fft_2048_16_5 is
port (
clock_c : in std_logic;
i1 : in  unsigned(0 downto 0);
i2 : in  unsigned(31 downto 0);
i3 : in  unsigned(31 downto 0);
i4 : in  unsigned(0 downto 0);
i5 : in  unsigned(0 downto 0);
o1 : out unsigned(0 downto 0);
o2 : out unsigned(31 downto 0);
o3 : out unsigned(31 downto 0));
end component cf_fft_2048_16_5;
component cf_fft_2048_16_2 is
port (
clock_c : in std_logic;
i1 : in  unsigned(0 downto 0);
i2 : in  unsigned(31 downto 0);
i3 : in  unsigned(31 downto 0);
i4 : in  unsigned(0 downto 0);
i5 : in  unsigned(0 downto 0);
o1 : out unsigned(0 downto 0);
o2 : out unsigned(31 downto 0);
o3 : out unsigned(31 downto 0));
end component cf_fft_2048_16_2;
begin
s1 : cf_fft_2048_16_25 port map (clock_c, s3_1, s3_2, s3_3, i4, i5, s1_1, s1_2, s1_3);
s2 : cf_fft_2048_16_8 port map (clock_c, s1_1, s1_2, s1_3, i4, i5, s2_1, s2_2, s2_3);
s3 : cf_fft_2048_16_6 port map (clock_c, s4_1, s4_2, s4_3, i4, i5, s3_1, s3_2, s3_3);
s4 : cf_fft_2048_16_5 port map (clock_c, s5_1, s5_2, s5_3, i4, i5, s4_1, s4_2, s4_3);
s5 : cf_fft_2048_16_2 port map (clock_c, i1, i2, i3, i4, i5, s5_1, s5_2, s5_3);
o3 <= s2_3;
o2 <= s2_2;
o1 <= s2_1;
end architecture rtl;

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
entity cf_fft_2048_16 is
port(
signal clock_c : in std_logic;
signal enable_i : in unsigned(0 downto 0);
signal reset_i : in unsigned(0 downto 0);
signal sync_i : in unsigned(0 downto 0);
signal data_0_i : in unsigned(31 downto 0);
signal data_1_i : in unsigned(31 downto 0);
signal sync_o : out unsigned(0 downto 0);
signal data_0_o : out unsigned(31 downto 0);
signal data_1_o : out unsigned(31 downto 0));
end entity cf_fft_2048_16;
architecture rtl of cf_fft_2048_16 is
component cf_fft_2048_16_1 is
port (
clock_c : in std_logic;
i1 : in  unsigned(0 downto 0);
i2 : in  unsigned(31 downto 0);
i3 : in  unsigned(31 downto 0);
i4 : in  unsigned(0 downto 0);
i5 : in  unsigned(0 downto 0);
o1 : out unsigned(0 downto 0);
o2 : out unsigned(31 downto 0);
o3 : out unsigned(31 downto 0));
end component cf_fft_2048_16_1;
signal n1 : unsigned(0 downto 0);
signal n2 : unsigned(31 downto 0);
signal n3 : unsigned(31 downto 0);
begin
s1 : cf_fft_2048_16_1 port map (clock_c, sync_i, data_0_i, data_1_i, enable_i, reset_i, n1, n2, n3);
sync_o <= n1;
data_0_o <= n2;
data_1_o <= n3;
end architecture rtl;


