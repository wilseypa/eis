--
--  Copyright (c) 2003 Launchbird Design Systems, Inc.
--  All rights reserved.
--  
--  Redistribution and use in source and binary forms, with or without modification, are permitted provided that the following conditions are met:
--    Redistributions of source code must retain the above copyright notice, this list of conditions and the following disclaimer.
--    Redistributions in binary form must reproduce the above copyright notice, this list of conditions and the following disclaimer in the documentation and/or other materials provided with the distribution.
--  
--  THIS SOFTWARE IS PROVIDED BY THE COPYRIGHT HOLDERS AND CONTRIBUTORS "AS IS" AND ANY EXPRESS OR IMPLIED WARRANTIES,
--  INCLUDING, BUT NOT LIMITED TO, THE IMPLIED WARRANTIES OF MERCHANTABILITY AND FITNESS FOR A PARTICULAR PURPOSE ARE DISCLAIMED.
--  IN NO EVENT SHALL THE COPYRIGHT OWNER OR CONTRIBUTORS BE LIABLE FOR ANY DIRECT, INDIRECT, INCIDENTAL, SPECIAL, EXEMPLARY,
--  OR CONSEQUENTIAL DAMAGES (INCLUDING, BUT NOT LIMITED TO, PROCUREMENT OF SUBSTITUTE GOODS OR SERVICES; LOSS OF USE, DATA, OR PROFITS;
--  OR BUSINESS INTERRUPTION) HOWEVER CAUSED AND ON ANY THEORY OF LIABILITY, WHETHER IN CONTRACT, STRICT LIABILITY, OR TORT
--  (INCLUDING NEGLIGENCE OR OTHERWISE) ARISING IN ANY WAY OUT OF THE USE OF THIS SOFTWARE, EVEN IF ADVISED OF THE POSSIBILITY OF SUCH DAMAGE.
--  
--  
--  Overview:
--  
--    Performs a radix 2 Fast Fourier Transform.
--    The FFT architecture is pipelined on a rank basis; each rank has its own butterfly and ranks are
--    isolated from each other using memory interleavers.  This FFT can perform calcualations on continuous
--    streaming data (one data set right after another).  More over, inputs and outputs are passed in pairs,
--    doubling the bandwidth.  For instance, a 2048 point FFT can perform a transform every 1024 cycles.
--  
--  Interface:
--  
--    Synchronization:
--      clock_c  : Clock input.
--      enable_i : Synchronous enable.
--      reset_i  : Synchronous reset.
--  
--    Inputs:
--      sync_i     : Input sync pulse must occur one frame prior to data input.
--      data_0_i   : Input data 0.  Width is 2 * precision.  Real on the left, imag on the right.
--      data_1_i   : Input data 1.  Width is 2 * precision.  Real on the left, imag on the right.
--  
--    Outputs:
--      sync_o     : Output sync pulse occurs one frame before data output.
--      data_0_o   : Output data 0.  Width is 2 * precision.  Real on the left, imag on the right.
--      data_1_o   : Output data 1.  Width is 2 * precision.  Real on the left, imag on the right.
--  
--  Built In Parameters:
--  
--    FFT Points   = 2048
--    Precision    = 8
--  
--  
--  
--  
--  Generated by Confluence 0.6.3  --  Launchbird Design Systems, Inc.  --  www.launchbird.com
--  
--  Build Date : Fri Aug 22 08:42:11 CDT 2003
--  
--  Interface
--  
--    Build Name    : cf_fft_2048_8
--    Clock Domains : clock_c  
--    Vector Input  : enable_i(1)
--    Vector Input  : reset_i(1)
--    Vector Input  : sync_i(1)
--    Vector Input  : data_0_i(16)
--    Vector Input  : data_1_i(16)
--    Vector Output : sync_o(1)
--    Vector Output : data_0_o(16)
--    Vector Output : data_1_o(16)
--  
--  
--  

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
entity cf_fft_2048_8_41 is
port (
clock_c : in std_logic;
i1 : in  unsigned(15 downto 0);
i2 : in  unsigned(15 downto 0);
i3 : in  unsigned(1 downto 0);
i4 : in  unsigned(0 downto 0);
i5 : in  unsigned(0 downto 0);
o1 : out unsigned(15 downto 0);
o2 : out unsigned(15 downto 0));
end entity cf_fft_2048_8_41;
architecture rtl of cf_fft_2048_8_41 is
signal n1 : unsigned(15 downto 0) := "0000000000000000";
signal n2 : unsigned(7 downto 0);
signal n3 : unsigned(7 downto 0);
signal n4 : unsigned(15 downto 0) := "0000000000000000";
signal n5 : unsigned(7 downto 0);
signal n6 : unsigned(7 downto 0);
signal n7 : unsigned(7 downto 0) := "00000000";
signal n8 : unsigned(7 downto 0) := "00000000";
signal n9 : unsigned(7 downto 0) := "00000000";
signal n10 : unsigned(7 downto 0) := "00000000";
signal n11 : unsigned(15 downto 0) := "0000000000000000";
signal n12 : unsigned(7 downto 0);
signal n13 : unsigned(7 downto 0);
signal n14 : unsigned(15 downto 0);
signal n15 : unsigned(7 downto 0);
signal n16 : unsigned(7 downto 0) := "00000000";
signal n17 : unsigned(15 downto 0);
signal n18 : unsigned(7 downto 0);
signal n19 : unsigned(7 downto 0) := "00000000";
signal n20 : unsigned(7 downto 0);
signal n21 : unsigned(7 downto 0) := "00000000";
signal n22 : unsigned(15 downto 0);
signal n23 : unsigned(7 downto 0);
signal n24 : unsigned(7 downto 0) := "00000000";
signal n25 : unsigned(15 downto 0);
signal n26 : unsigned(7 downto 0);
signal n27 : unsigned(7 downto 0) := "00000000";
signal n28 : unsigned(7 downto 0);
signal n29 : unsigned(7 downto 0) := "00000000";
signal n30 : unsigned(7 downto 0);
signal n31 : unsigned(7 downto 0);
signal n32 : unsigned(15 downto 0);
signal n33 : unsigned(15 downto 0) := "0000000000000000";
signal n34 : unsigned(7 downto 0);
signal n35 : unsigned(7 downto 0);
signal n36 : unsigned(15 downto 0);
signal n37 : unsigned(15 downto 0) := "0000000000000000";
begin
process (clock_c) begin
  if rising_edge(clock_c) then
    if i5 = "1" then
      n1 <= "0000000000000000";
    elsif i4 = "1" then
      n1 <= i1;
    end if;
  end if;
end process;
n2 <= n1(15 downto 15) &
  n1(14 downto 14) &
  n1(13 downto 13) &
  n1(12 downto 12) &
  n1(11 downto 11) &
  n1(10 downto 10) &
  n1(9 downto 9) &
  n1(8 downto 8);
n3 <= n1(7 downto 7) &
  n1(6 downto 6) &
  n1(5 downto 5) &
  n1(4 downto 4) &
  n1(3 downto 3) &
  n1(2 downto 2) &
  n1(1 downto 1) &
  n1(0 downto 0);
process (clock_c) begin
  if rising_edge(clock_c) then
    if i5 = "1" then
      n4 <= "0000000000000000";
    elsif i4 = "1" then
      n4 <= i2;
    end if;
  end if;
end process;
n5 <= n4(15 downto 15) &
  n4(14 downto 14) &
  n4(13 downto 13) &
  n4(12 downto 12) &
  n4(11 downto 11) &
  n4(10 downto 10) &
  n4(9 downto 9) &
  n4(8 downto 8);
n6 <= n4(7 downto 7) &
  n4(6 downto 6) &
  n4(5 downto 5) &
  n4(4 downto 4) &
  n4(3 downto 3) &
  n4(2 downto 2) &
  n4(1 downto 1) &
  n4(0 downto 0);
process (clock_c) begin
  if rising_edge(clock_c) then
    if i5 = "1" then
      n7 <= "00000000";
    elsif i4 = "1" then
      n7 <= n2;
    end if;
  end if;
end process;
process (clock_c) begin
  if rising_edge(clock_c) then
    if i5 = "1" then
      n8 <= "00000000";
    elsif i4 = "1" then
      n8 <= n7;
    end if;
  end if;
end process;
process (clock_c) begin
  if rising_edge(clock_c) then
    if i5 = "1" then
      n9 <= "00000000";
    elsif i4 = "1" then
      n9 <= n3;
    end if;
  end if;
end process;
process (clock_c) begin
  if rising_edge(clock_c) then
    if i5 = "1" then
      n10 <= "00000000";
    elsif i4 = "1" then
      n10 <= n9;
    end if;
  end if;
end process;
process (clock_c) begin
  if rising_edge(clock_c) then 
    if i4 = "1" then
      case i3 is
        when "00" => n11 <= "0111111100000000";
        when "01" => n11 <= "0101101010100101";
        when "10" => n11 <= "0000000010000000";
        when "11" => n11 <= "1010010110100101";
        when others => n11 <= "XXXXXXXXXXXXXXXX";
      end case;
    end if;
  end if;
end process;
n12 <= n11(15 downto 15) &
  n11(14 downto 14) &
  n11(13 downto 13) &
  n11(12 downto 12) &
  n11(11 downto 11) &
  n11(10 downto 10) &
  n11(9 downto 9) &
  n11(8 downto 8);
n13 <= n11(7 downto 7) &
  n11(6 downto 6) &
  n11(5 downto 5) &
  n11(4 downto 4) &
  n11(3 downto 3) &
  n11(2 downto 2) &
  n11(1 downto 1) &
  n11(0 downto 0);
n14 <= unsigned(signed(n5) * signed(n12));
n15 <= n14(14 downto 14) &
  n14(13 downto 13) &
  n14(12 downto 12) &
  n14(11 downto 11) &
  n14(10 downto 10) &
  n14(9 downto 9) &
  n14(8 downto 8) &
  n14(7 downto 7);
process (clock_c) begin
  if rising_edge(clock_c) then
    if i5 = "1" then
      n16 <= "00000000";
    elsif i4 = "1" then
      n16 <= n15;
    end if;
  end if;
end process;
n17 <= unsigned(signed(n6) * signed(n13));
n18 <= n17(14 downto 14) &
  n17(13 downto 13) &
  n17(12 downto 12) &
  n17(11 downto 11) &
  n17(10 downto 10) &
  n17(9 downto 9) &
  n17(8 downto 8) &
  n17(7 downto 7);
process (clock_c) begin
  if rising_edge(clock_c) then
    if i5 = "1" then
      n19 <= "00000000";
    elsif i4 = "1" then
      n19 <= n18;
    end if;
  end if;
end process;
n20 <= n16 - n19;
process (clock_c) begin
  if rising_edge(clock_c) then
    if i5 = "1" then
      n21 <= "00000000";
    elsif i4 = "1" then
      n21 <= n20;
    end if;
  end if;
end process;
n22 <= unsigned(signed(n5) * signed(n13));
n23 <= n22(14 downto 14) &
  n22(13 downto 13) &
  n22(12 downto 12) &
  n22(11 downto 11) &
  n22(10 downto 10) &
  n22(9 downto 9) &
  n22(8 downto 8) &
  n22(7 downto 7);
process (clock_c) begin
  if rising_edge(clock_c) then
    if i5 = "1" then
      n24 <= "00000000";
    elsif i4 = "1" then
      n24 <= n23;
    end if;
  end if;
end process;
n25 <= unsigned(signed(n6) * signed(n12));
n26 <= n25(14 downto 14) &
  n25(13 downto 13) &
  n25(12 downto 12) &
  n25(11 downto 11) &
  n25(10 downto 10) &
  n25(9 downto 9) &
  n25(8 downto 8) &
  n25(7 downto 7);
process (clock_c) begin
  if rising_edge(clock_c) then
    if i5 = "1" then
      n27 <= "00000000";
    elsif i4 = "1" then
      n27 <= n26;
    end if;
  end if;
end process;
n28 <= n24 + n27;
process (clock_c) begin
  if rising_edge(clock_c) then
    if i5 = "1" then
      n29 <= "00000000";
    elsif i4 = "1" then
      n29 <= n28;
    end if;
  end if;
end process;
n30 <= n8 + n21;
n31 <= n10 + n29;
n32 <= n30 & n31;
process (clock_c) begin
  if rising_edge(clock_c) then
    if i5 = "1" then
      n33 <= "0000000000000000";
    elsif i4 = "1" then
      n33 <= n32;
    end if;
  end if;
end process;
n34 <= n8 - n21;
n35 <= n10 - n29;
n36 <= n34 & n35;
process (clock_c) begin
  if rising_edge(clock_c) then
    if i5 = "1" then
      n37 <= "0000000000000000";
    elsif i4 = "1" then
      n37 <= n36;
    end if;
  end if;
end process;
o2 <= n37;
o1 <= n33;
end architecture rtl;

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
entity cf_fft_2048_8_40 is
port (
i1 : in  unsigned(0 downto 0);
i2 : in  unsigned(0 downto 0);
i3 : in  unsigned(0 downto 0);
i4 : in  unsigned(0 downto 0);
i5 : in  unsigned(2 downto 0);
o1 : out unsigned(0 downto 0));
end entity cf_fft_2048_8_40;
architecture rtl of cf_fft_2048_8_40 is
signal n1 : unsigned(2 downto 0);
signal n2 : unsigned(2 downto 0);
signal n3 : unsigned(2 downto 0);
signal n4 : unsigned(0 downto 0);
signal n5 : unsigned(0 downto 0);
signal n6 : unsigned(0 downto 0);
signal n7 : unsigned(0 downto 0);
signal n8 : unsigned(0 downto 0);
signal n9 : unsigned(0 downto 0);
begin
n1 <= "001";
n2 <= "011";
n3 <= "101";
n4 <= "1" when i5 = n1 else "0";
n5 <= "1" when i5 = n2 else "0";
n6 <= "1" when i5 = n3 else "0";
n7 <= i2 when n6 = "1" else i1;
n8 <= i3 when n5 = "1" else n7;
n9 <= i4 when n4 = "1" else n8;
o1 <= n9;
end architecture rtl;

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
entity cf_fft_2048_8_39 is
port (
i1 : in  unsigned(0 downto 0);
i2 : in  unsigned(0 downto 0);
i3 : in  unsigned(0 downto 0);
i4 : in  unsigned(0 downto 0);
i5 : in  unsigned(0 downto 0);
i6 : in  unsigned(0 downto 0);
i7 : in  unsigned(0 downto 0);
i8 : in  unsigned(2 downto 0);
o1 : out unsigned(0 downto 0));
end entity cf_fft_2048_8_39;
architecture rtl of cf_fft_2048_8_39 is
signal n1 : unsigned(2 downto 0);
signal n2 : unsigned(2 downto 0);
signal n3 : unsigned(2 downto 0);
signal n4 : unsigned(0 downto 0);
signal n5 : unsigned(0 downto 0);
signal n6 : unsigned(0 downto 0);
signal n7 : unsigned(0 downto 0);
signal n8 : unsigned(0 downto 0);
signal n9 : unsigned(0 downto 0);
signal s10_1 : unsigned(0 downto 0);
component cf_fft_2048_8_40 is
port (
i1 : in  unsigned(0 downto 0);
i2 : in  unsigned(0 downto 0);
i3 : in  unsigned(0 downto 0);
i4 : in  unsigned(0 downto 0);
i5 : in  unsigned(2 downto 0);
o1 : out unsigned(0 downto 0));
end component cf_fft_2048_8_40;
begin
n1 <= "010";
n2 <= "100";
n3 <= "110";
n4 <= "1" when i8 = n1 else "0";
n5 <= "1" when i8 = n2 else "0";
n6 <= "1" when i8 = n3 else "0";
n7 <= i5 when n6 = "1" else s10_1;
n8 <= i6 when n5 = "1" else n7;
n9 <= i7 when n4 = "1" else n8;
s10 : cf_fft_2048_8_40 port map (i1, i2, i3, i4, i8, s10_1);
o1 <= n9;
end architecture rtl;

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
entity cf_fft_2048_8_38 is
port (
o1 : out unsigned(0 downto 0);
o2 : out unsigned(0 downto 0);
o3 : out unsigned(0 downto 0);
o4 : out unsigned(0 downto 0);
o5 : out unsigned(0 downto 0);
o6 : out unsigned(0 downto 0);
o7 : out unsigned(0 downto 0);
o8 : out unsigned(0 downto 0));
end entity cf_fft_2048_8_38;
architecture rtl of cf_fft_2048_8_38 is
signal n1 : unsigned(0 downto 0);
signal n2 : unsigned(0 downto 0);
signal n3 : unsigned(0 downto 0);
signal n4 : unsigned(0 downto 0);
signal n5 : unsigned(0 downto 0);
signal n6 : unsigned(0 downto 0);
signal n7 : unsigned(0 downto 0);
signal n8 : unsigned(0 downto 0);
begin
n1 <= "0";
n2 <= "1";
n3 <= "0";
n4 <= "1";
n5 <= "0";
n6 <= "1";
n7 <= "0";
n8 <= "0";
o8 <= n8;
o7 <= n7;
o6 <= n6;
o5 <= n5;
o4 <= n4;
o3 <= n3;
o2 <= n2;
o1 <= n1;
end architecture rtl;

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
entity cf_fft_2048_8_37 is
port (
i1 : in  unsigned(0 downto 0);
i2 : in  unsigned(0 downto 0);
i3 : in  unsigned(0 downto 0);
i4 : in  unsigned(2 downto 0);
o1 : out unsigned(0 downto 0));
end entity cf_fft_2048_8_37;
architecture rtl of cf_fft_2048_8_37 is
signal n1 : unsigned(2 downto 0);
signal n2 : unsigned(2 downto 0);
signal n3 : unsigned(2 downto 0);
signal n4 : unsigned(0 downto 0);
signal n5 : unsigned(0 downto 0);
signal n6 : unsigned(0 downto 0);
signal n7 : unsigned(0 downto 0);
signal n8 : unsigned(0 downto 0);
signal n9 : unsigned(0 downto 0);
signal n10 : unsigned(0 downto 0);
begin
n1 <= "010";
n2 <= "100";
n3 <= "110";
n4 <= "1" when i4 = n1 else "0";
n5 <= "1" when i4 = n2 else "0";
n6 <= "1" when i4 = n3 else "0";
n7 <= i1 when n6 = "1" else n10;
n8 <= i2 when n5 = "1" else n7;
n9 <= i3 when n4 = "1" else n8;
n10 <= "1";
o1 <= n9;
end architecture rtl;

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
entity cf_fft_2048_8_36 is
port (
i1 : in  unsigned(2 downto 0);
o1 : out unsigned(0 downto 0));
end entity cf_fft_2048_8_36;
architecture rtl of cf_fft_2048_8_36 is
signal n1 : unsigned(0 downto 0);
signal n2 : unsigned(0 downto 0);
signal n3 : unsigned(0 downto 0);
signal n4 : unsigned(0 downto 0);
signal n5 : unsigned(2 downto 0);
signal n6 : unsigned(0 downto 0);
signal n7 : unsigned(0 downto 0);
signal s8_1 : unsigned(0 downto 0);
component cf_fft_2048_8_37 is
port (
i1 : in  unsigned(0 downto 0);
i2 : in  unsigned(0 downto 0);
i3 : in  unsigned(0 downto 0);
i4 : in  unsigned(2 downto 0);
o1 : out unsigned(0 downto 0));
end component cf_fft_2048_8_37;
begin
n1 <= "0";
n2 <= "0";
n3 <= "0";
n4 <= "0";
n5 <= "000";
n6 <= "1" when i1 = n5 else "0";
n7 <= n4 when n6 = "1" else s8_1;
s8 : cf_fft_2048_8_37 port map (n1, n2, n3, i1, s8_1);
o1 <= n7;
end architecture rtl;

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
entity cf_fft_2048_8_35 is
port (
clock_c : in std_logic;
i1 : in  unsigned(1 downto 0);
i2 : in  unsigned(0 downto 0);
i3 : in  unsigned(0 downto 0);
o1 : out unsigned(0 downto 0));
end entity cf_fft_2048_8_35;
architecture rtl of cf_fft_2048_8_35 is
signal n1 : unsigned(2 downto 0);
signal n2 : unsigned(2 downto 0);
signal n3 : unsigned(0 downto 0);
signal n4 : unsigned(0 downto 0);
signal n5 : unsigned(0 downto 0) := "0";
signal s6_1 : unsigned(0 downto 0);
signal s7_1 : unsigned(0 downto 0);
signal s7_2 : unsigned(0 downto 0);
signal s7_3 : unsigned(0 downto 0);
signal s7_4 : unsigned(0 downto 0);
signal s7_5 : unsigned(0 downto 0);
signal s7_6 : unsigned(0 downto 0);
signal s7_7 : unsigned(0 downto 0);
signal s7_8 : unsigned(0 downto 0);
signal s8_1 : unsigned(0 downto 0);
component cf_fft_2048_8_39 is
port (
i1 : in  unsigned(0 downto 0);
i2 : in  unsigned(0 downto 0);
i3 : in  unsigned(0 downto 0);
i4 : in  unsigned(0 downto 0);
i5 : in  unsigned(0 downto 0);
i6 : in  unsigned(0 downto 0);
i7 : in  unsigned(0 downto 0);
i8 : in  unsigned(2 downto 0);
o1 : out unsigned(0 downto 0));
end component cf_fft_2048_8_39;
component cf_fft_2048_8_38 is
port (
o1 : out unsigned(0 downto 0);
o2 : out unsigned(0 downto 0);
o3 : out unsigned(0 downto 0);
o4 : out unsigned(0 downto 0);
o5 : out unsigned(0 downto 0);
o6 : out unsigned(0 downto 0);
o7 : out unsigned(0 downto 0);
o8 : out unsigned(0 downto 0));
end component cf_fft_2048_8_38;
component cf_fft_2048_8_36 is
port (
i1 : in  unsigned(2 downto 0);
o1 : out unsigned(0 downto 0));
end component cf_fft_2048_8_36;
begin
n1 <= "000";
n2 <= i1 & n5;
n3 <= "1" when n2 = n1 else "0";
n4 <= s7_8 when n3 = "1" else s6_1;
process (clock_c) begin
  if rising_edge(clock_c) then
    if i3 = "1" then
      n5 <= "0";
    elsif i2 = "1" then
      n5 <= n4;
    end if;
  end if;
end process;
s6 : cf_fft_2048_8_39 port map (s7_1, s7_2, s7_3, s7_4, s7_5, s7_6, s7_7, n2, s6_1);
s7 : cf_fft_2048_8_38 port map (s7_1, s7_2, s7_3, s7_4, s7_5, s7_6, s7_7, s7_8);
s8 : cf_fft_2048_8_36 port map (n2, s8_1);
o1 <= s8_1;
end architecture rtl;

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
entity cf_fft_2048_8_34 is
port (
i1 : in  unsigned(0 downto 0);
i2 : in  unsigned(0 downto 0);
i3 : in  unsigned(0 downto 0);
i4 : in  unsigned(0 downto 0);
i5 : in  unsigned(1 downto 0);
o1 : out unsigned(0 downto 0));
end entity cf_fft_2048_8_34;
architecture rtl of cf_fft_2048_8_34 is
signal n1 : unsigned(1 downto 0);
signal n2 : unsigned(1 downto 0);
signal n3 : unsigned(1 downto 0);
signal n4 : unsigned(0 downto 0);
signal n5 : unsigned(0 downto 0);
signal n6 : unsigned(0 downto 0);
signal n7 : unsigned(0 downto 0);
signal n8 : unsigned(0 downto 0);
signal n9 : unsigned(0 downto 0);
begin
n1 <= "00";
n2 <= "10";
n3 <= "01";
n4 <= "1" when i5 = n1 else "0";
n5 <= "1" when i5 = n2 else "0";
n6 <= "1" when i5 = n3 else "0";
n7 <= i2 when n6 = "1" else i1;
n8 <= i3 when n5 = "1" else n7;
n9 <= i4 when n4 = "1" else n8;
o1 <= n9;
end architecture rtl;

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
entity cf_fft_2048_8_33 is
port (
i1 : in  unsigned(1 downto 0);
o1 : out unsigned(0 downto 0));
end entity cf_fft_2048_8_33;
architecture rtl of cf_fft_2048_8_33 is
signal n1 : unsigned(0 downto 0);
signal n2 : unsigned(0 downto 0);
signal n3 : unsigned(1 downto 0);
signal n4 : unsigned(1 downto 0);
signal n5 : unsigned(0 downto 0);
signal n6 : unsigned(0 downto 0);
signal n7 : unsigned(0 downto 0);
signal n8 : unsigned(0 downto 0);
signal n9 : unsigned(0 downto 0);
begin
n1 <= "0";
n2 <= "0";
n3 <= "00";
n4 <= "10";
n5 <= "1" when i1 = n3 else "0";
n6 <= "1" when i1 = n4 else "0";
n7 <= n1 when n6 = "1" else n9;
n8 <= n2 when n5 = "1" else n7;
n9 <= "1";
o1 <= n8;
end architecture rtl;

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
entity cf_fft_2048_8_32 is
port (
clock_c : in std_logic;
i1 : in  unsigned(0 downto 0);
i2 : in  unsigned(0 downto 0);
i3 : in  unsigned(0 downto 0);
o1 : out unsigned(0 downto 0));
end entity cf_fft_2048_8_32;
architecture rtl of cf_fft_2048_8_32 is
signal n1 : unsigned(0 downto 0);
signal n2 : unsigned(0 downto 0);
signal n3 : unsigned(0 downto 0);
signal n4 : unsigned(0 downto 0);
signal n5 : unsigned(1 downto 0);
signal n6 : unsigned(0 downto 0) := "0";
signal s7_1 : unsigned(0 downto 0);
signal s8_1 : unsigned(0 downto 0);
component cf_fft_2048_8_34 is
port (
i1 : in  unsigned(0 downto 0);
i2 : in  unsigned(0 downto 0);
i3 : in  unsigned(0 downto 0);
i4 : in  unsigned(0 downto 0);
i5 : in  unsigned(1 downto 0);
o1 : out unsigned(0 downto 0));
end component cf_fft_2048_8_34;
component cf_fft_2048_8_33 is
port (
i1 : in  unsigned(1 downto 0);
o1 : out unsigned(0 downto 0));
end component cf_fft_2048_8_33;
begin
n1 <= "0";
n2 <= "1";
n3 <= "1";
n4 <= "0";
n5 <= i1 & n6;
process (clock_c) begin
  if rising_edge(clock_c) then
    if i3 = "1" then
      n6 <= "0";
    elsif i2 = "1" then
      n6 <= s7_1;
    end if;
  end if;
end process;
s7 : cf_fft_2048_8_34 port map (n1, n2, n3, n4, n5, s7_1);
s8 : cf_fft_2048_8_33 port map (n5, s8_1);
o1 <= s8_1;
end architecture rtl;

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
entity cf_fft_2048_8_31 is
port (
clock_c : in std_logic;
i1 : in  unsigned(31 downto 0);
i2 : in  unsigned(0 downto 0);
i3 : in  unsigned(8 downto 0);
i4 : in  unsigned(0 downto 0);
i5 : in  unsigned(0 downto 0);
i6 : in  unsigned(0 downto 0);
o1 : out unsigned(31 downto 0));
end entity cf_fft_2048_8_31;
architecture rtl of cf_fft_2048_8_31 is
signal n1 : unsigned(8 downto 0);
signal n2 : unsigned(8 downto 0);
signal n3 : unsigned(8 downto 0) := "000000000";
signal n4 : unsigned(0 downto 0);
signal n5 : unsigned(0 downto 0);
signal n6 : unsigned(31 downto 0);
signal n6a : unsigned(8 downto 0) := "000000000";
type   n6mt is array (511 downto 0) of unsigned(31 downto 0);
signal n6m : n6mt;
signal n7 : unsigned(0 downto 0);
signal n8 : unsigned(31 downto 0);
signal n8a : unsigned(8 downto 0) := "000000000";
type   n8mt is array (511 downto 0) of unsigned(31 downto 0);
signal n8m : n8mt;
signal n9 : unsigned(0 downto 0) := "0";
signal n10 : unsigned(31 downto 0);
signal n11 : unsigned(0 downto 0);
signal s12_1 : unsigned(0 downto 0);
component cf_fft_2048_8_32 is
port (
clock_c : in std_logic;
i1 : in  unsigned(0 downto 0);
i2 : in  unsigned(0 downto 0);
i3 : in  unsigned(0 downto 0);
o1 : out unsigned(0 downto 0));
end component cf_fft_2048_8_32;
begin
n1 <= "000000001";
n2 <= n3 + n1;
process (clock_c) begin
  if rising_edge(clock_c) then
    if n11 = "1" then
      n3 <= "000000000";
    elsif i5 = "1" then
      n3 <= n2;
    end if;
  end if;
end process;
n4 <= not s12_1;
n5 <= i4 and n4;
process (clock_c) begin
  if rising_edge(clock_c) then
    if i5 = "1" then
      if n5 = "1" then
        n6m(to_integer(i3)) <= i1;
      end if;
      n6a <= n3;
    end if;
  end if;
end process;
n6 <= n6m(to_integer(n6a));
n7 <= i4 and s12_1;
process (clock_c) begin
  if rising_edge(clock_c) then
    if i5 = "1" then
      if n7 = "1" then
        n8m(to_integer(i3)) <= i1;
      end if;
      n8a <= n3;
    end if;
  end if;
end process;
n8 <= n8m(to_integer(n8a));
process (clock_c) begin
  if rising_edge(clock_c) then
    if i6 = "1" then
      n9 <= "0";
    elsif i5 = "1" then
      n9 <= n4;
    end if;
  end if;
end process;
n10 <= n8 when n9 = "1" else n6;
n11 <= i2 or i6;
s12 : cf_fft_2048_8_32 port map (clock_c, i2, i5, i6, s12_1);
o1 <= n10;
end architecture rtl;

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
entity cf_fft_2048_8_30 is
port (
clock_c : in std_logic;
i1 : in  unsigned(31 downto 0);
i2 : in  unsigned(0 downto 0);
i3 : in  unsigned(8 downto 0);
i4 : in  unsigned(0 downto 0);
i5 : in  unsigned(0 downto 0);
i6 : in  unsigned(0 downto 0);
o1 : out unsigned(0 downto 0);
o2 : out unsigned(0 downto 0);
o3 : out unsigned(31 downto 0));
end entity cf_fft_2048_8_30;
architecture rtl of cf_fft_2048_8_30 is
signal n1 : unsigned(8 downto 0);
signal n2 : unsigned(8 downto 0);
signal n3 : unsigned(8 downto 0) := "000000000";
signal n4 : unsigned(0 downto 0);
signal n5 : unsigned(0 downto 0) := "0";
signal n6 : unsigned(8 downto 0);
signal n7 : unsigned(0 downto 0);
signal n8 : unsigned(0 downto 0);
signal n9 : unsigned(31 downto 0);
signal n9a : unsigned(8 downto 0) := "000000000";
type   n9mt is array (511 downto 0) of unsigned(31 downto 0);
signal n9m : n9mt;
signal n10 : unsigned(0 downto 0);
signal n11 : unsigned(31 downto 0);
signal n11a : unsigned(8 downto 0) := "000000000";
type   n11mt is array (511 downto 0) of unsigned(31 downto 0);
signal n11m : n11mt;
signal n12 : unsigned(0 downto 0) := "0";
signal n13 : unsigned(31 downto 0);
signal n14 : unsigned(0 downto 0);
signal s15_1 : unsigned(0 downto 0);
component cf_fft_2048_8_32 is
port (
clock_c : in std_logic;
i1 : in  unsigned(0 downto 0);
i2 : in  unsigned(0 downto 0);
i3 : in  unsigned(0 downto 0);
o1 : out unsigned(0 downto 0));
end component cf_fft_2048_8_32;
begin
n1 <= "000000001";
n2 <= n3 + n1;
process (clock_c) begin
  if rising_edge(clock_c) then
    if n14 = "1" then
      n3 <= "000000000";
    elsif i5 = "1" then
      n3 <= n2;
    end if;
  end if;
end process;
n4 <= not s15_1;
process (clock_c) begin
  if rising_edge(clock_c) then
    if i6 = "1" then
      n5 <= "0";
    elsif i5 = "1" then
      n5 <= i2;
    end if;
  end if;
end process;
n6 <= "000000000";
n7 <= "1" when n3 = n6 else "0";
n8 <= i4 and n4;
process (clock_c) begin
  if rising_edge(clock_c) then
    if i5 = "1" then
      if n8 = "1" then
        n9m(to_integer(i3)) <= i1;
      end if;
      n9a <= n3;
    end if;
  end if;
end process;
n9 <= n9m(to_integer(n9a));
n10 <= i4 and s15_1;
process (clock_c) begin
  if rising_edge(clock_c) then
    if i5 = "1" then
      if n10 = "1" then
        n11m(to_integer(i3)) <= i1;
      end if;
      n11a <= n3;
    end if;
  end if;
end process;
n11 <= n11m(to_integer(n11a));
process (clock_c) begin
  if rising_edge(clock_c) then
    if i6 = "1" then
      n12 <= "0";
    elsif i5 = "1" then
      n12 <= n4;
    end if;
  end if;
end process;
n13 <= n11 when n12 = "1" else n9;
n14 <= i2 or i6;
s15 : cf_fft_2048_8_32 port map (clock_c, i2, i5, i6, s15_1);
o3 <= n13;
o2 <= n7;
o1 <= n5;
end architecture rtl;

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
entity cf_fft_2048_8_29 is
port (
i1 : in  unsigned(0 downto 0);
i2 : in  unsigned(0 downto 0);
i3 : in  unsigned(0 downto 0);
i4 : in  unsigned(2 downto 0);
o1 : out unsigned(0 downto 0));
end entity cf_fft_2048_8_29;
architecture rtl of cf_fft_2048_8_29 is
signal n1 : unsigned(2 downto 0);
signal n2 : unsigned(2 downto 0);
signal n3 : unsigned(2 downto 0);
signal n4 : unsigned(0 downto 0);
signal n5 : unsigned(0 downto 0);
signal n6 : unsigned(0 downto 0);
signal n7 : unsigned(0 downto 0);
signal n8 : unsigned(0 downto 0);
signal n9 : unsigned(0 downto 0);
signal n10 : unsigned(0 downto 0);
begin
n1 <= "110";
n2 <= "001";
n3 <= "011";
n4 <= "1" when i4 = n1 else "0";
n5 <= "1" when i4 = n2 else "0";
n6 <= "1" when i4 = n3 else "0";
n7 <= i1 when n6 = "1" else n10;
n8 <= i2 when n5 = "1" else n7;
n9 <= i3 when n4 = "1" else n8;
n10 <= "1";
o1 <= n9;
end architecture rtl;

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
entity cf_fft_2048_8_28 is
port (
i1 : in  unsigned(0 downto 0);
i2 : in  unsigned(0 downto 0);
i3 : in  unsigned(0 downto 0);
i4 : in  unsigned(0 downto 0);
i5 : in  unsigned(0 downto 0);
i6 : in  unsigned(0 downto 0);
i7 : in  unsigned(2 downto 0);
o1 : out unsigned(0 downto 0));
end entity cf_fft_2048_8_28;
architecture rtl of cf_fft_2048_8_28 is
signal n1 : unsigned(2 downto 0);
signal n2 : unsigned(2 downto 0);
signal n3 : unsigned(2 downto 0);
signal n4 : unsigned(0 downto 0);
signal n5 : unsigned(0 downto 0);
signal n6 : unsigned(0 downto 0);
signal n7 : unsigned(0 downto 0);
signal n8 : unsigned(0 downto 0);
signal n9 : unsigned(0 downto 0);
signal s10_1 : unsigned(0 downto 0);
component cf_fft_2048_8_29 is
port (
i1 : in  unsigned(0 downto 0);
i2 : in  unsigned(0 downto 0);
i3 : in  unsigned(0 downto 0);
i4 : in  unsigned(2 downto 0);
o1 : out unsigned(0 downto 0));
end component cf_fft_2048_8_29;
begin
n1 <= "000";
n2 <= "010";
n3 <= "100";
n4 <= "1" when i7 = n1 else "0";
n5 <= "1" when i7 = n2 else "0";
n6 <= "1" when i7 = n3 else "0";
n7 <= i4 when n6 = "1" else s10_1;
n8 <= i5 when n5 = "1" else n7;
n9 <= i6 when n4 = "1" else n8;
s10 : cf_fft_2048_8_29 port map (i1, i2, i3, i7, s10_1);
o1 <= n9;
end architecture rtl;

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
entity cf_fft_2048_8_27 is
port (
clock_c : in std_logic;
i1 : in  unsigned(1 downto 0);
i2 : in  unsigned(0 downto 0);
i3 : in  unsigned(0 downto 0);
o1 : out unsigned(0 downto 0));
end entity cf_fft_2048_8_27;
architecture rtl of cf_fft_2048_8_27 is
signal n1 : unsigned(0 downto 0);
signal n2 : unsigned(0 downto 0);
signal n3 : unsigned(0 downto 0);
signal n4 : unsigned(0 downto 0);
signal n5 : unsigned(0 downto 0);
signal n6 : unsigned(0 downto 0);
signal n7 : unsigned(0 downto 0);
signal n8 : unsigned(0 downto 0);
signal n9 : unsigned(0 downto 0);
signal n10 : unsigned(0 downto 0);
signal n11 : unsigned(0 downto 0);
signal n12 : unsigned(0 downto 0);
signal n13 : unsigned(2 downto 0);
signal n14 : unsigned(0 downto 0) := "0";
signal s15_1 : unsigned(0 downto 0);
signal s16_1 : unsigned(0 downto 0);
component cf_fft_2048_8_28 is
port (
i1 : in  unsigned(0 downto 0);
i2 : in  unsigned(0 downto 0);
i3 : in  unsigned(0 downto 0);
i4 : in  unsigned(0 downto 0);
i5 : in  unsigned(0 downto 0);
i6 : in  unsigned(0 downto 0);
i7 : in  unsigned(2 downto 0);
o1 : out unsigned(0 downto 0));
end component cf_fft_2048_8_28;
begin
n1 <= "0";
n2 <= "1";
n3 <= "1";
n4 <= "1";
n5 <= "0";
n6 <= "0";
n7 <= "0";
n8 <= "1";
n9 <= "1";
n10 <= "1";
n11 <= "0";
n12 <= "0";
n13 <= i1 & n14;
process (clock_c) begin
  if rising_edge(clock_c) then
    if i3 = "1" then
      n14 <= "0";
    elsif i2 = "1" then
      n14 <= s15_1;
    end if;
  end if;
end process;
s15 : cf_fft_2048_8_28 port map (n1, n2, n3, n4, n5, n6, n13, s15_1);
s16 : cf_fft_2048_8_28 port map (n7, n8, n9, n10, n11, n12, n13, s16_1);
o1 <= s16_1;
end architecture rtl;

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
entity cf_fft_2048_8_26 is
port (
clock_c : in std_logic;
i1 : in  unsigned(0 downto 0);
i2 : in  unsigned(0 downto 0);
i3 : in  unsigned(0 downto 0);
o1 : out unsigned(9 downto 0);
o2 : out unsigned(0 downto 0));
end entity cf_fft_2048_8_26;
architecture rtl of cf_fft_2048_8_26 is
signal n1 : unsigned(9 downto 0);
signal n2 : unsigned(9 downto 0);
signal n3 : unsigned(9 downto 0) := "0000000000";
signal n4 : unsigned(9 downto 0);
signal n5 : unsigned(0 downto 0);
signal n6 : unsigned(1 downto 0);
signal n7 : unsigned(0 downto 0) := "0";
signal n8 : unsigned(0 downto 0);
signal n9 : unsigned(0 downto 0);
signal n10 : unsigned(0 downto 0);
signal s11_1 : unsigned(0 downto 0);
component cf_fft_2048_8_27 is
port (
clock_c : in std_logic;
i1 : in  unsigned(1 downto 0);
i2 : in  unsigned(0 downto 0);
i3 : in  unsigned(0 downto 0);
o1 : out unsigned(0 downto 0));
end component cf_fft_2048_8_27;
begin
n1 <= "0000000001";
n2 <= n3 + n1;
process (clock_c) begin
  if rising_edge(clock_c) then
    if n9 = "1" then
      n3 <= "0000000000";
    elsif n10 = "1" then
      n3 <= n2;
    end if;
  end if;
end process;
n4 <= "1111111111";
n5 <= "1" when n3 = n4 else "0";
n6 <= i1 & n5;
process (clock_c) begin
  if rising_edge(clock_c) then
    if i3 = "1" then
      n7 <= "0";
    elsif i2 = "1" then
      n7 <= s11_1;
    end if;
  end if;
end process;
n8 <= n7 and n5;
n9 <= i1 or i3;
n10 <= s11_1 and i2;
s11 : cf_fft_2048_8_27 port map (clock_c, n6, i2, i3, s11_1);
o2 <= n8;
o1 <= n3;
end architecture rtl;

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
entity cf_fft_2048_8_25 is
port (
clock_c : in std_logic;
i1 : in  unsigned(0 downto 0);
i2 : in  unsigned(15 downto 0);
i3 : in  unsigned(15 downto 0);
i4 : in  unsigned(0 downto 0);
i5 : in  unsigned(0 downto 0);
o1 : out unsigned(0 downto 0);
o2 : out unsigned(15 downto 0);
o3 : out unsigned(15 downto 0));
end entity cf_fft_2048_8_25;
architecture rtl of cf_fft_2048_8_25 is
signal n1 : unsigned(1 downto 0);
signal n2 : unsigned(31 downto 0);
signal n3 : unsigned(0 downto 0) := "0";
signal n4 : unsigned(0 downto 0) := "0";
signal n5 : unsigned(0 downto 0) := "0";
signal n6 : unsigned(0 downto 0) := "0";
signal n7 : unsigned(8 downto 0);
signal n8 : unsigned(8 downto 0) := "000000000";
signal n9 : unsigned(8 downto 0) := "000000000";
signal n10 : unsigned(8 downto 0) := "000000000";
signal n11 : unsigned(8 downto 0) := "000000000";
signal n12 : unsigned(0 downto 0);
signal n13 : unsigned(0 downto 0) := "0";
signal n14 : unsigned(0 downto 0) := "0";
signal n15 : unsigned(0 downto 0) := "0";
signal n16 : unsigned(0 downto 0) := "0";
signal n17 : unsigned(0 downto 0);
signal n18 : unsigned(1 downto 0);
signal n19 : unsigned(15 downto 0);
signal n20 : unsigned(15 downto 0);
signal n21 : unsigned(15 downto 0);
signal n22 : unsigned(15 downto 0);
signal n23 : unsigned(15 downto 0);
signal n24 : unsigned(15 downto 0);
signal s25_1 : unsigned(15 downto 0);
signal s25_2 : unsigned(15 downto 0);
signal s26_1 : unsigned(0 downto 0);
signal s27_1 : unsigned(31 downto 0);
signal s28_1 : unsigned(0 downto 0);
signal s28_2 : unsigned(0 downto 0);
signal s28_3 : unsigned(31 downto 0);
signal s29_1 : unsigned(9 downto 0);
signal s29_2 : unsigned(0 downto 0);
component cf_fft_2048_8_41 is
port (
clock_c : in std_logic;
i1 : in  unsigned(15 downto 0);
i2 : in  unsigned(15 downto 0);
i3 : in  unsigned(1 downto 0);
i4 : in  unsigned(0 downto 0);
i5 : in  unsigned(0 downto 0);
o1 : out unsigned(15 downto 0);
o2 : out unsigned(15 downto 0));
end component cf_fft_2048_8_41;
component cf_fft_2048_8_35 is
port (
clock_c : in std_logic;
i1 : in  unsigned(1 downto 0);
i2 : in  unsigned(0 downto 0);
i3 : in  unsigned(0 downto 0);
o1 : out unsigned(0 downto 0));
end component cf_fft_2048_8_35;
component cf_fft_2048_8_31 is
port (
clock_c : in std_logic;
i1 : in  unsigned(31 downto 0);
i2 : in  unsigned(0 downto 0);
i3 : in  unsigned(8 downto 0);
i4 : in  unsigned(0 downto 0);
i5 : in  unsigned(0 downto 0);
i6 : in  unsigned(0 downto 0);
o1 : out unsigned(31 downto 0));
end component cf_fft_2048_8_31;
component cf_fft_2048_8_30 is
port (
clock_c : in std_logic;
i1 : in  unsigned(31 downto 0);
i2 : in  unsigned(0 downto 0);
i3 : in  unsigned(8 downto 0);
i4 : in  unsigned(0 downto 0);
i5 : in  unsigned(0 downto 0);
i6 : in  unsigned(0 downto 0);
o1 : out unsigned(0 downto 0);
o2 : out unsigned(0 downto 0);
o3 : out unsigned(31 downto 0));
end component cf_fft_2048_8_30;
component cf_fft_2048_8_26 is
port (
clock_c : in std_logic;
i1 : in  unsigned(0 downto 0);
i2 : in  unsigned(0 downto 0);
i3 : in  unsigned(0 downto 0);
o1 : out unsigned(9 downto 0);
o2 : out unsigned(0 downto 0));
end component cf_fft_2048_8_26;
begin
n1 <= s29_1(9 downto 9) &
  s29_1(8 downto 8);
n2 <= s25_1 & s25_2;
process (clock_c) begin
  if rising_edge(clock_c) then
    if i5 = "1" then
      n3 <= "0";
    elsif i4 = "1" then
      n3 <= s29_2;
    end if;
  end if;
end process;
process (clock_c) begin
  if rising_edge(clock_c) then
    if i5 = "1" then
      n4 <= "0";
    elsif i4 = "1" then
      n4 <= n3;
    end if;
  end if;
end process;
process (clock_c) begin
  if rising_edge(clock_c) then
    if i5 = "1" then
      n5 <= "0";
    elsif i4 = "1" then
      n5 <= n4;
    end if;
  end if;
end process;
process (clock_c) begin
  if rising_edge(clock_c) then
    if i5 = "1" then
      n6 <= "0";
    elsif i4 = "1" then
      n6 <= n5;
    end if;
  end if;
end process;
n7 <= s29_1(9 downto 9) &
  s29_1(8 downto 8) &
  s29_1(7 downto 7) &
  s29_1(6 downto 6) &
  s29_1(5 downto 5) &
  s29_1(4 downto 4) &
  s29_1(3 downto 3) &
  s29_1(2 downto 2) &
  s29_1(1 downto 1);
process (clock_c) begin
  if rising_edge(clock_c) then
    if i5 = "1" then
      n8 <= "000000000";
    elsif i4 = "1" then
      n8 <= n7;
    end if;
  end if;
end process;
process (clock_c) begin
  if rising_edge(clock_c) then
    if i5 = "1" then
      n9 <= "000000000";
    elsif i4 = "1" then
      n9 <= n8;
    end if;
  end if;
end process;
process (clock_c) begin
  if rising_edge(clock_c) then
    if i5 = "1" then
      n10 <= "000000000";
    elsif i4 = "1" then
      n10 <= n9;
    end if;
  end if;
end process;
process (clock_c) begin
  if rising_edge(clock_c) then
    if i5 = "1" then
      n11 <= "000000000";
    elsif i4 = "1" then
      n11 <= n10;
    end if;
  end if;
end process;
n12 <= s29_1(0 downto 0);
process (clock_c) begin
  if rising_edge(clock_c) then
    if i5 = "1" then
      n13 <= "0";
    elsif i4 = "1" then
      n13 <= n12;
    end if;
  end if;
end process;
process (clock_c) begin
  if rising_edge(clock_c) then
    if i5 = "1" then
      n14 <= "0";
    elsif i4 = "1" then
      n14 <= n13;
    end if;
  end if;
end process;
process (clock_c) begin
  if rising_edge(clock_c) then
    if i5 = "1" then
      n15 <= "0";
    elsif i4 = "1" then
      n15 <= n14;
    end if;
  end if;
end process;
process (clock_c) begin
  if rising_edge(clock_c) then
    if i5 = "1" then
      n16 <= "0";
    elsif i4 = "1" then
      n16 <= n15;
    end if;
  end if;
end process;
n17 <= not n16;
n18 <= s28_2 & s28_1;
n19 <= s28_3(31 downto 31) &
  s28_3(30 downto 30) &
  s28_3(29 downto 29) &
  s28_3(28 downto 28) &
  s28_3(27 downto 27) &
  s28_3(26 downto 26) &
  s28_3(25 downto 25) &
  s28_3(24 downto 24) &
  s28_3(23 downto 23) &
  s28_3(22 downto 22) &
  s28_3(21 downto 21) &
  s28_3(20 downto 20) &
  s28_3(19 downto 19) &
  s28_3(18 downto 18) &
  s28_3(17 downto 17) &
  s28_3(16 downto 16);
n20 <= s28_3(15 downto 15) &
  s28_3(14 downto 14) &
  s28_3(13 downto 13) &
  s28_3(12 downto 12) &
  s28_3(11 downto 11) &
  s28_3(10 downto 10) &
  s28_3(9 downto 9) &
  s28_3(8 downto 8) &
  s28_3(7 downto 7) &
  s28_3(6 downto 6) &
  s28_3(5 downto 5) &
  s28_3(4 downto 4) &
  s28_3(3 downto 3) &
  s28_3(2 downto 2) &
  s28_3(1 downto 1) &
  s28_3(0 downto 0);
n21 <= s27_1(31 downto 31) &
  s27_1(30 downto 30) &
  s27_1(29 downto 29) &
  s27_1(28 downto 28) &
  s27_1(27 downto 27) &
  s27_1(26 downto 26) &
  s27_1(25 downto 25) &
  s27_1(24 downto 24) &
  s27_1(23 downto 23) &
  s27_1(22 downto 22) &
  s27_1(21 downto 21) &
  s27_1(20 downto 20) &
  s27_1(19 downto 19) &
  s27_1(18 downto 18) &
  s27_1(17 downto 17) &
  s27_1(16 downto 16);
n22 <= s27_1(15 downto 15) &
  s27_1(14 downto 14) &
  s27_1(13 downto 13) &
  s27_1(12 downto 12) &
  s27_1(11 downto 11) &
  s27_1(10 downto 10) &
  s27_1(9 downto 9) &
  s27_1(8 downto 8) &
  s27_1(7 downto 7) &
  s27_1(6 downto 6) &
  s27_1(5 downto 5) &
  s27_1(4 downto 4) &
  s27_1(3 downto 3) &
  s27_1(2 downto 2) &
  s27_1(1 downto 1) &
  s27_1(0 downto 0);
n23 <= n20 when s26_1 = "1" else n19;
n24 <= n22 when s26_1 = "1" else n21;
s25 : cf_fft_2048_8_41 port map (clock_c, i2, i3, n1, i4, i5, s25_1, s25_2);
s26 : cf_fft_2048_8_35 port map (clock_c, n18, i4, i5, s26_1);
s27 : cf_fft_2048_8_31 port map (clock_c, n2, n6, n11, n16, i4, i5, s27_1);
s28 : cf_fft_2048_8_30 port map (clock_c, n2, n6, n11, n17, i4, i5, s28_1, s28_2, s28_3);
s29 : cf_fft_2048_8_26 port map (clock_c, i1, i4, i5, s29_1, s29_2);
o3 <= n24;
o2 <= n23;
o1 <= s28_1;
end architecture rtl;

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
entity cf_fft_2048_8_24 is
port (
clock_c : in std_logic;
i1 : in  unsigned(15 downto 0);
i2 : in  unsigned(15 downto 0);
i3 : in  unsigned(9 downto 0);
i4 : in  unsigned(0 downto 0);
i5 : in  unsigned(0 downto 0);
o1 : out unsigned(15 downto 0);
o2 : out unsigned(15 downto 0));
end entity cf_fft_2048_8_24;
architecture rtl of cf_fft_2048_8_24 is
signal n1 : unsigned(15 downto 0) := "0000000000000000";
signal n2 : unsigned(7 downto 0);
signal n3 : unsigned(7 downto 0);
signal n4 : unsigned(15 downto 0) := "0000000000000000";
signal n5 : unsigned(7 downto 0);
signal n6 : unsigned(7 downto 0);
signal n7 : unsigned(7 downto 0) := "00000000";
signal n8 : unsigned(7 downto 0) := "00000000";
signal n9 : unsigned(7 downto 0) := "00000000";
signal n10 : unsigned(7 downto 0) := "00000000";
signal n11 : unsigned(15 downto 0) := "0000000000000000";
signal n12 : unsigned(7 downto 0);
signal n13 : unsigned(7 downto 0);
signal n14 : unsigned(15 downto 0);
signal n15 : unsigned(7 downto 0);
signal n16 : unsigned(7 downto 0) := "00000000";
signal n17 : unsigned(15 downto 0);
signal n18 : unsigned(7 downto 0);
signal n19 : unsigned(7 downto 0) := "00000000";
signal n20 : unsigned(7 downto 0);
signal n21 : unsigned(7 downto 0) := "00000000";
signal n22 : unsigned(15 downto 0);
signal n23 : unsigned(7 downto 0);
signal n24 : unsigned(7 downto 0) := "00000000";
signal n25 : unsigned(15 downto 0);
signal n26 : unsigned(7 downto 0);
signal n27 : unsigned(7 downto 0) := "00000000";
signal n28 : unsigned(7 downto 0);
signal n29 : unsigned(7 downto 0) := "00000000";
signal n30 : unsigned(7 downto 0);
signal n31 : unsigned(7 downto 0);
signal n32 : unsigned(15 downto 0);
signal n33 : unsigned(15 downto 0) := "0000000000000000";
signal n34 : unsigned(7 downto 0);
signal n35 : unsigned(7 downto 0);
signal n36 : unsigned(15 downto 0);
signal n37 : unsigned(15 downto 0) := "0000000000000000";
begin
process (clock_c) begin
  if rising_edge(clock_c) then
    if i5 = "1" then
      n1 <= "0000000000000000";
    elsif i4 = "1" then
      n1 <= i1;
    end if;
  end if;
end process;
n2 <= n1(15 downto 15) &
  n1(14 downto 14) &
  n1(13 downto 13) &
  n1(12 downto 12) &
  n1(11 downto 11) &
  n1(10 downto 10) &
  n1(9 downto 9) &
  n1(8 downto 8);
n3 <= n1(7 downto 7) &
  n1(6 downto 6) &
  n1(5 downto 5) &
  n1(4 downto 4) &
  n1(3 downto 3) &
  n1(2 downto 2) &
  n1(1 downto 1) &
  n1(0 downto 0);
process (clock_c) begin
  if rising_edge(clock_c) then
    if i5 = "1" then
      n4 <= "0000000000000000";
    elsif i4 = "1" then
      n4 <= i2;
    end if;
  end if;
end process;
n5 <= n4(15 downto 15) &
  n4(14 downto 14) &
  n4(13 downto 13) &
  n4(12 downto 12) &
  n4(11 downto 11) &
  n4(10 downto 10) &
  n4(9 downto 9) &
  n4(8 downto 8);
n6 <= n4(7 downto 7) &
  n4(6 downto 6) &
  n4(5 downto 5) &
  n4(4 downto 4) &
  n4(3 downto 3) &
  n4(2 downto 2) &
  n4(1 downto 1) &
  n4(0 downto 0);
process (clock_c) begin
  if rising_edge(clock_c) then
    if i5 = "1" then
      n7 <= "00000000";
    elsif i4 = "1" then
      n7 <= n2;
    end if;
  end if;
end process;
process (clock_c) begin
  if rising_edge(clock_c) then
    if i5 = "1" then
      n8 <= "00000000";
    elsif i4 = "1" then
      n8 <= n7;
    end if;
  end if;
end process;
process (clock_c) begin
  if rising_edge(clock_c) then
    if i5 = "1" then
      n9 <= "00000000";
    elsif i4 = "1" then
      n9 <= n3;
    end if;
  end if;
end process;
process (clock_c) begin
  if rising_edge(clock_c) then
    if i5 = "1" then
      n10 <= "00000000";
    elsif i4 = "1" then
      n10 <= n9;
    end if;
  end if;
end process;
process (clock_c) begin
  if rising_edge(clock_c) then 
    if i4 = "1" then
      case i3 is
        when "0000000000" => n11 <= "0111111100000000";
        when "0000000001" => n11 <= "0111111111111111";
        when "0000000010" => n11 <= "0111111111111111";
        when "0000000011" => n11 <= "0111111111111110";
        when "0000000100" => n11 <= "0111111111111110";
        when "0000000101" => n11 <= "0111111111111110";
        when "0000000110" => n11 <= "0111111111111101";
        when "0000000111" => n11 <= "0111111111111101";
        when "0000001000" => n11 <= "0111111111111100";
        when "0000001001" => n11 <= "0111111111111100";
        when "0000001010" => n11 <= "0111111111111100";
        when "0000001011" => n11 <= "0111111111111011";
        when "0000001100" => n11 <= "0111111111111011";
        when "0000001101" => n11 <= "0111111111111010";
        when "0000001110" => n11 <= "0111111111111010";
        when "0000001111" => n11 <= "0111111111111010";
        when "0000010000" => n11 <= "0111111111111001";
        when "0000010001" => n11 <= "0111111111111001";
        when "0000010010" => n11 <= "0111111111111000";
        when "0000010011" => n11 <= "0111111111111000";
        when "0000010100" => n11 <= "0111111111111000";
        when "0000010101" => n11 <= "0111111111110111";
        when "0000010110" => n11 <= "0111111111110111";
        when "0000010111" => n11 <= "0111111111110110";
        when "0000011000" => n11 <= "0111111111110110";
        when "0000011001" => n11 <= "0111111111110110";
        when "0000011010" => n11 <= "0111111111110101";
        when "0000011011" => n11 <= "0111111111110101";
        when "0000011100" => n11 <= "0111111111110101";
        when "0000011101" => n11 <= "0111111111110100";
        when "0000011110" => n11 <= "0111111111110100";
        when "0000011111" => n11 <= "0111111111110011";
        when "0000100000" => n11 <= "0111111111110011";
        when "0000100001" => n11 <= "0111111111110011";
        when "0000100010" => n11 <= "0111111111110010";
        when "0000100011" => n11 <= "0111111111110010";
        when "0000100100" => n11 <= "0111111111110001";
        when "0000100101" => n11 <= "0111111111110001";
        when "0000100110" => n11 <= "0111111111110001";
        when "0000100111" => n11 <= "0111111111110000";
        when "0000101000" => n11 <= "0111111111110000";
        when "0000101001" => n11 <= "0111111011101111";
        when "0000101010" => n11 <= "0111111011101111";
        when "0000101011" => n11 <= "0111111011101111";
        when "0000101100" => n11 <= "0111111011101110";
        when "0000101101" => n11 <= "0111111011101110";
        when "0000101110" => n11 <= "0111111011101101";
        when "0000101111" => n11 <= "0111111011101101";
        when "0000110000" => n11 <= "0111111011101101";
        when "0000110001" => n11 <= "0111111011101100";
        when "0000110010" => n11 <= "0111111011101100";
        when "0000110011" => n11 <= "0111111011101100";
        when "0000110100" => n11 <= "0111111011101011";
        when "0000110101" => n11 <= "0111111011101011";
        when "0000110110" => n11 <= "0111111011101010";
        when "0000110111" => n11 <= "0111111011101010";
        when "0000111000" => n11 <= "0111111011101010";
        when "0000111001" => n11 <= "0111111011101001";
        when "0000111010" => n11 <= "0111110111101001";
        when "0000111011" => n11 <= "0111110111101000";
        when "0000111100" => n11 <= "0111110111101000";
        when "0000111101" => n11 <= "0111110111101000";
        when "0000111110" => n11 <= "0111110111100111";
        when "0000111111" => n11 <= "0111110111100111";
        when "0001000000" => n11 <= "0111110111100111";
        when "0001000001" => n11 <= "0111110111100110";
        when "0001000010" => n11 <= "0111110111100110";
        when "0001000011" => n11 <= "0111110111100101";
        when "0001000100" => n11 <= "0111110111100101";
        when "0001000101" => n11 <= "0111110111100101";
        when "0001000110" => n11 <= "0111110111100100";
        when "0001000111" => n11 <= "0111110011100100";
        when "0001001000" => n11 <= "0111110011100011";
        when "0001001001" => n11 <= "0111110011100011";
        when "0001001010" => n11 <= "0111110011100011";
        when "0001001011" => n11 <= "0111110011100010";
        when "0001001100" => n11 <= "0111110011100010";
        when "0001001101" => n11 <= "0111110011100010";
        when "0001001110" => n11 <= "0111110011100001";
        when "0001001111" => n11 <= "0111110011100001";
        when "0001010000" => n11 <= "0111110011100000";
        when "0001010001" => n11 <= "0111110011100000";
        when "0001010010" => n11 <= "0111101111100000";
        when "0001010011" => n11 <= "0111101111011111";
        when "0001010100" => n11 <= "0111101111011111";
        when "0001010101" => n11 <= "0111101111011110";
        when "0001010110" => n11 <= "0111101111011110";
        when "0001010111" => n11 <= "0111101111011110";
        when "0001011000" => n11 <= "0111101111011101";
        when "0001011001" => n11 <= "0111101111011101";
        when "0001011010" => n11 <= "0111101111011101";
        when "0001011011" => n11 <= "0111101111011100";
        when "0001011100" => n11 <= "0111101011011100";
        when "0001011101" => n11 <= "0111101011011011";
        when "0001011110" => n11 <= "0111101011011011";
        when "0001011111" => n11 <= "0111101011011011";
        when "0001100000" => n11 <= "0111101011011010";
        when "0001100001" => n11 <= "0111101011011010";
        when "0001100010" => n11 <= "0111101011011010";
        when "0001100011" => n11 <= "0111101011011001";
        when "0001100100" => n11 <= "0111101011011001";
        when "0001100101" => n11 <= "0111100111011000";
        when "0001100110" => n11 <= "0111100111011000";
        when "0001100111" => n11 <= "0111100111011000";
        when "0001101000" => n11 <= "0111100111010111";
        when "0001101001" => n11 <= "0111100111010111";
        when "0001101010" => n11 <= "0111100111010111";
        when "0001101011" => n11 <= "0111100111010110";
        when "0001101100" => n11 <= "0111100111010110";
        when "0001101101" => n11 <= "0111100011010101";
        when "0001101110" => n11 <= "0111100011010101";
        when "0001101111" => n11 <= "0111100011010101";
        when "0001110000" => n11 <= "0111100011010100";
        when "0001110001" => n11 <= "0111100011010100";
        when "0001110010" => n11 <= "0111100011010100";
        when "0001110011" => n11 <= "0111100011010011";
        when "0001110100" => n11 <= "0111011111010011";
        when "0001110101" => n11 <= "0111011111010011";
        when "0001110110" => n11 <= "0111011111010010";
        when "0001110111" => n11 <= "0111011111010010";
        when "0001111000" => n11 <= "0111011111010001";
        when "0001111001" => n11 <= "0111011111010001";
        when "0001111010" => n11 <= "0111011111010001";
        when "0001111011" => n11 <= "0111011011010000";
        when "0001111100" => n11 <= "0111011011010000";
        when "0001111101" => n11 <= "0111011011010000";
        when "0001111110" => n11 <= "0111011011001111";
        when "0001111111" => n11 <= "0111011011001111";
        when "0010000000" => n11 <= "0111011011001111";
        when "0010000001" => n11 <= "0111011011001110";
        when "0010000010" => n11 <= "0111010111001110";
        when "0010000011" => n11 <= "0111010111001101";
        when "0010000100" => n11 <= "0111010111001101";
        when "0010000101" => n11 <= "0111010111001101";
        when "0010000110" => n11 <= "0111010111001100";
        when "0010000111" => n11 <= "0111010111001100";
        when "0010001000" => n11 <= "0111010111001100";
        when "0010001001" => n11 <= "0111010011001011";
        when "0010001010" => n11 <= "0111010011001011";
        when "0010001011" => n11 <= "0111010011001011";
        when "0010001100" => n11 <= "0111010011001010";
        when "0010001101" => n11 <= "0111010011001010";
        when "0010001110" => n11 <= "0111010011001001";
        when "0010001111" => n11 <= "0111001111001001";
        when "0010010000" => n11 <= "0111001111001001";
        when "0010010001" => n11 <= "0111001111001000";
        when "0010010010" => n11 <= "0111001111001000";
        when "0010010011" => n11 <= "0111001111001000";
        when "0010010100" => n11 <= "0111001111000111";
        when "0010010101" => n11 <= "0111001011000111";
        when "0010010110" => n11 <= "0111001011000111";
        when "0010010111" => n11 <= "0111001011000110";
        when "0010011000" => n11 <= "0111001011000110";
        when "0010011001" => n11 <= "0111001011000110";
        when "0010011010" => n11 <= "0111000111000101";
        when "0010011011" => n11 <= "0111000111000101";
        when "0010011100" => n11 <= "0111000111000101";
        when "0010011101" => n11 <= "0111000111000100";
        when "0010011110" => n11 <= "0111000111000100";
        when "0010011111" => n11 <= "0111000111000100";
        when "0010100000" => n11 <= "0111000011000011";
        when "0010100001" => n11 <= "0111000011000011";
        when "0010100010" => n11 <= "0111000011000010";
        when "0010100011" => n11 <= "0111000011000010";
        when "0010100100" => n11 <= "0111000011000010";
        when "0010100101" => n11 <= "0110111111000001";
        when "0010100110" => n11 <= "0110111111000001";
        when "0010100111" => n11 <= "0110111111000001";
        when "0010101000" => n11 <= "0110111111000000";
        when "0010101001" => n11 <= "0110111111000000";
        when "0010101010" => n11 <= "0110111011000000";
        when "0010101011" => n11 <= "0110111010111111";
        when "0010101100" => n11 <= "0110111010111111";
        when "0010101101" => n11 <= "0110111010111111";
        when "0010101110" => n11 <= "0110111010111110";
        when "0010101111" => n11 <= "0110110110111110";
        when "0010110000" => n11 <= "0110110110111110";
        when "0010110001" => n11 <= "0110110110111101";
        when "0010110010" => n11 <= "0110110110111101";
        when "0010110011" => n11 <= "0110110110111101";
        when "0010110100" => n11 <= "0110110010111100";
        when "0010110101" => n11 <= "0110110010111100";
        when "0010110110" => n11 <= "0110110010111100";
        when "0010110111" => n11 <= "0110110010111011";
        when "0010111000" => n11 <= "0110110010111011";
        when "0010111001" => n11 <= "0110101110111011";
        when "0010111010" => n11 <= "0110101110111010";
        when "0010111011" => n11 <= "0110101110111010";
        when "0010111100" => n11 <= "0110101110111010";
        when "0010111101" => n11 <= "0110101110111001";
        when "0010111110" => n11 <= "0110101010111001";
        when "0010111111" => n11 <= "0110101010111001";
        when "0011000000" => n11 <= "0110101010111000";
        when "0011000001" => n11 <= "0110101010111000";
        when "0011000010" => n11 <= "0110100110111000";
        when "0011000011" => n11 <= "0110100110110111";
        when "0011000100" => n11 <= "0110100110110111";
        when "0011000101" => n11 <= "0110100110110111";
        when "0011000110" => n11 <= "0110100110110110";
        when "0011000111" => n11 <= "0110100010110110";
        when "0011001000" => n11 <= "0110100010110110";
        when "0011001001" => n11 <= "0110100010110101";
        when "0011001010" => n11 <= "0110100010110101";
        when "0011001011" => n11 <= "0110011110110101";
        when "0011001100" => n11 <= "0110011110110101";
        when "0011001101" => n11 <= "0110011110110100";
        when "0011001110" => n11 <= "0110011110110100";
        when "0011001111" => n11 <= "0110011110110100";
        when "0011010000" => n11 <= "0110011010110011";
        when "0011010001" => n11 <= "0110011010110011";
        when "0011010010" => n11 <= "0110011010110011";
        when "0011010011" => n11 <= "0110011010110010";
        when "0011010100" => n11 <= "0110010110110010";
        when "0011010101" => n11 <= "0110010110110010";
        when "0011010110" => n11 <= "0110010110110001";
        when "0011010111" => n11 <= "0110010110110001";
        when "0011011000" => n11 <= "0110010010110001";
        when "0011011001" => n11 <= "0110010010110000";
        when "0011011010" => n11 <= "0110010010110000";
        when "0011011011" => n11 <= "0110010010110000";
        when "0011011100" => n11 <= "0110001110110000";
        when "0011011101" => n11 <= "0110001110101111";
        when "0011011110" => n11 <= "0110001110101111";
        when "0011011111" => n11 <= "0110001110101111";
        when "0011100000" => n11 <= "0110001010101110";
        when "0011100001" => n11 <= "0110001010101110";
        when "0011100010" => n11 <= "0110001010101110";
        when "0011100011" => n11 <= "0110001010101101";
        when "0011100100" => n11 <= "0110000110101101";
        when "0011100101" => n11 <= "0110000110101101";
        when "0011100110" => n11 <= "0110000110101100";
        when "0011100111" => n11 <= "0110000110101100";
        when "0011101000" => n11 <= "0110000010101100";
        when "0011101001" => n11 <= "0110000010101100";
        when "0011101010" => n11 <= "0110000010101011";
        when "0011101011" => n11 <= "0110000010101011";
        when "0011101100" => n11 <= "0101111110101011";
        when "0011101101" => n11 <= "0101111110101010";
        when "0011101110" => n11 <= "0101111110101010";
        when "0011101111" => n11 <= "0101111110101010";
        when "0011110000" => n11 <= "0101111010101010";
        when "0011110001" => n11 <= "0101111010101001";
        when "0011110010" => n11 <= "0101111010101001";
        when "0011110011" => n11 <= "0101111010101001";
        when "0011110100" => n11 <= "0101110110101000";
        when "0011110101" => n11 <= "0101110110101000";
        when "0011110110" => n11 <= "0101110110101000";
        when "0011110111" => n11 <= "0101110010101000";
        when "0011111000" => n11 <= "0101110010100111";
        when "0011111001" => n11 <= "0101110010100111";
        when "0011111010" => n11 <= "0101110010100111";
        when "0011111011" => n11 <= "0101101110100110";
        when "0011111100" => n11 <= "0101101110100110";
        when "0011111101" => n11 <= "0101101110100110";
        when "0011111110" => n11 <= "0101101110100110";
        when "0011111111" => n11 <= "0101101010100101";
        when "0100000000" => n11 <= "0101101010100101";
        when "0100000001" => n11 <= "0101101010100101";
        when "0100000010" => n11 <= "0101100110100100";
        when "0100000011" => n11 <= "0101100110100100";
        when "0100000100" => n11 <= "0101100110100100";
        when "0100000101" => n11 <= "0101100110100100";
        when "0100000110" => n11 <= "0101100010100011";
        when "0100000111" => n11 <= "0101100010100011";
        when "0100001000" => n11 <= "0101100010100011";
        when "0100001001" => n11 <= "0101011110100011";
        when "0100001010" => n11 <= "0101011110100010";
        when "0100001011" => n11 <= "0101011110100010";
        when "0100001100" => n11 <= "0101011110100010";
        when "0100001101" => n11 <= "0101011010100001";
        when "0100001110" => n11 <= "0101011010100001";
        when "0100001111" => n11 <= "0101011010100001";
        when "0100010000" => n11 <= "0101010110100001";
        when "0100010001" => n11 <= "0101010110100000";
        when "0100010010" => n11 <= "0101010110100000";
        when "0100010011" => n11 <= "0101010110100000";
        when "0100010100" => n11 <= "0101010010100000";
        when "0100010101" => n11 <= "0101010010011111";
        when "0100010110" => n11 <= "0101010010011111";
        when "0100010111" => n11 <= "0101001110011111";
        when "0100011000" => n11 <= "0101001110011111";
        when "0100011001" => n11 <= "0101001110011110";
        when "0100011010" => n11 <= "0101001110011110";
        when "0100011011" => n11 <= "0101001010011110";
        when "0100011100" => n11 <= "0101001010011110";
        when "0100011101" => n11 <= "0101001010011101";
        when "0100011110" => n11 <= "0101000110011101";
        when "0100011111" => n11 <= "0101000110011101";
        when "0100100000" => n11 <= "0101000110011101";
        when "0100100001" => n11 <= "0101000010011100";
        when "0100100010" => n11 <= "0101000010011100";
        when "0100100011" => n11 <= "0101000010011100";
        when "0100100100" => n11 <= "0100111110011100";
        when "0100100101" => n11 <= "0100111110011011";
        when "0100100110" => n11 <= "0100111110011011";
        when "0100100111" => n11 <= "0100111110011011";
        when "0100101000" => n11 <= "0100111010011011";
        when "0100101001" => n11 <= "0100111010011010";
        when "0100101010" => n11 <= "0100111010011010";
        when "0100101011" => n11 <= "0100110110011010";
        when "0100101100" => n11 <= "0100110110011010";
        when "0100101101" => n11 <= "0100110110011001";
        when "0100101110" => n11 <= "0100110010011001";
        when "0100101111" => n11 <= "0100110010011001";
        when "0100110000" => n11 <= "0100110010011001";
        when "0100110001" => n11 <= "0100101110011000";
        when "0100110010" => n11 <= "0100101110011000";
        when "0100110011" => n11 <= "0100101110011000";
        when "0100110100" => n11 <= "0100101010011000";
        when "0100110101" => n11 <= "0100101010011000";
        when "0100110110" => n11 <= "0100101010010111";
        when "0100110111" => n11 <= "0100101010010111";
        when "0100111000" => n11 <= "0100100110010111";
        when "0100111001" => n11 <= "0100100110010111";
        when "0100111010" => n11 <= "0100100110010110";
        when "0100111011" => n11 <= "0100100010010110";
        when "0100111100" => n11 <= "0100100010010110";
        when "0100111101" => n11 <= "0100100010010110";
        when "0100111110" => n11 <= "0100011110010110";
        when "0100111111" => n11 <= "0100011110010101";
        when "0101000000" => n11 <= "0100011110010101";
        when "0101000001" => n11 <= "0100011010010101";
        when "0101000010" => n11 <= "0100011010010101";
        when "0101000011" => n11 <= "0100011010010100";
        when "0101000100" => n11 <= "0100010110010100";
        when "0101000101" => n11 <= "0100010110010100";
        when "0101000110" => n11 <= "0100010110010100";
        when "0101000111" => n11 <= "0100010010010100";
        when "0101001000" => n11 <= "0100010010010011";
        when "0101001001" => n11 <= "0100010010010011";
        when "0101001010" => n11 <= "0100001110010011";
        when "0101001011" => n11 <= "0100001110010011";
        when "0101001100" => n11 <= "0100001110010011";
        when "0101001101" => n11 <= "0100001010010010";
        when "0101001110" => n11 <= "0100001010010010";
        when "0101001111" => n11 <= "0100001010010010";
        when "0101010000" => n11 <= "0100000110010010";
        when "0101010001" => n11 <= "0100000110010010";
        when "0101010010" => n11 <= "0100000110010001";
        when "0101010011" => n11 <= "0100000010010001";
        when "0101010100" => n11 <= "0100000010010001";
        when "0101010101" => n11 <= "0100000010010001";
        when "0101010110" => n11 <= "0011111110010001";
        when "0101010111" => n11 <= "0011111110010000";
        when "0101011000" => n11 <= "0011111110010000";
        when "0101011001" => n11 <= "0011111010010000";
        when "0101011010" => n11 <= "0011111010010000";
        when "0101011011" => n11 <= "0011111010010000";
        when "0101011100" => n11 <= "0011110110001111";
        when "0101011101" => n11 <= "0011110110001111";
        when "0101011110" => n11 <= "0011110110001111";
        when "0101011111" => n11 <= "0011110010001111";
        when "0101100000" => n11 <= "0011110010001111";
        when "0101100001" => n11 <= "0011101110001110";
        when "0101100010" => n11 <= "0011101110001110";
        when "0101100011" => n11 <= "0011101110001110";
        when "0101100100" => n11 <= "0011101010001110";
        when "0101100101" => n11 <= "0011101010001110";
        when "0101100110" => n11 <= "0011101010001110";
        when "0101100111" => n11 <= "0011100110001101";
        when "0101101000" => n11 <= "0011100110001101";
        when "0101101001" => n11 <= "0011100110001101";
        when "0101101010" => n11 <= "0011100010001101";
        when "0101101011" => n11 <= "0011100010001101";
        when "0101101100" => n11 <= "0011100010001100";
        when "0101101101" => n11 <= "0011011110001100";
        when "0101101110" => n11 <= "0011011110001100";
        when "0101101111" => n11 <= "0011011110001100";
        when "0101110000" => n11 <= "0011011010001100";
        when "0101110001" => n11 <= "0011011010001100";
        when "0101110010" => n11 <= "0011011010001011";
        when "0101110011" => n11 <= "0011010110001011";
        when "0101110100" => n11 <= "0011010110001011";
        when "0101110101" => n11 <= "0011010010001011";
        when "0101110110" => n11 <= "0011010010001011";
        when "0101110111" => n11 <= "0011010010001011";
        when "0101111000" => n11 <= "0011001110001010";
        when "0101111001" => n11 <= "0011001110001010";
        when "0101111010" => n11 <= "0011001110001010";
        when "0101111011" => n11 <= "0011001010001010";
        when "0101111100" => n11 <= "0011001010001010";
        when "0101111101" => n11 <= "0011001010001010";
        when "0101111110" => n11 <= "0011000110001010";
        when "0101111111" => n11 <= "0011000110001001";
        when "0110000000" => n11 <= "0011000010001001";
        when "0110000001" => n11 <= "0011000010001001";
        when "0110000010" => n11 <= "0011000010001001";
        when "0110000011" => n11 <= "0010111110001001";
        when "0110000100" => n11 <= "0010111110001001";
        when "0110000101" => n11 <= "0010111110001001";
        when "0110000110" => n11 <= "0010111010001000";
        when "0110000111" => n11 <= "0010111010001000";
        when "0110001000" => n11 <= "0010111010001000";
        when "0110001001" => n11 <= "0010110110001000";
        when "0110001010" => n11 <= "0010110110001000";
        when "0110001011" => n11 <= "0010110010001000";
        when "0110001100" => n11 <= "0010110010001000";
        when "0110001101" => n11 <= "0010110010000111";
        when "0110001110" => n11 <= "0010101110000111";
        when "0110001111" => n11 <= "0010101110000111";
        when "0110010000" => n11 <= "0010101110000111";
        when "0110010001" => n11 <= "0010101010000111";
        when "0110010010" => n11 <= "0010101010000111";
        when "0110010011" => n11 <= "0010101010000111";
        when "0110010100" => n11 <= "0010100110000110";
        when "0110010101" => n11 <= "0010100110000110";
        when "0110010110" => n11 <= "0010100010000110";
        when "0110010111" => n11 <= "0010100010000110";
        when "0110011000" => n11 <= "0010100010000110";
        when "0110011001" => n11 <= "0010011110000110";
        when "0110011010" => n11 <= "0010011110000110";
        when "0110011011" => n11 <= "0010011110000110";
        when "0110011100" => n11 <= "0010011010000101";
        when "0110011101" => n11 <= "0010011010000101";
        when "0110011110" => n11 <= "0010010110000101";
        when "0110011111" => n11 <= "0010010110000101";
        when "0110100000" => n11 <= "0010010110000101";
        when "0110100001" => n11 <= "0010010010000101";
        when "0110100010" => n11 <= "0010010010000101";
        when "0110100011" => n11 <= "0010010010000101";
        when "0110100100" => n11 <= "0010001110000101";
        when "0110100101" => n11 <= "0010001110000100";
        when "0110100110" => n11 <= "0010001010000100";
        when "0110100111" => n11 <= "0010001010000100";
        when "0110101000" => n11 <= "0010001010000100";
        when "0110101001" => n11 <= "0010000110000100";
        when "0110101010" => n11 <= "0010000110000100";
        when "0110101011" => n11 <= "0010000110000100";
        when "0110101100" => n11 <= "0010000010000100";
        when "0110101101" => n11 <= "0010000010000100";
        when "0110101110" => n11 <= "0001111110000100";
        when "0110101111" => n11 <= "0001111110000011";
        when "0110110000" => n11 <= "0001111110000011";
        when "0110110001" => n11 <= "0001111010000011";
        when "0110110010" => n11 <= "0001111010000011";
        when "0110110011" => n11 <= "0001110110000011";
        when "0110110100" => n11 <= "0001110110000011";
        when "0110110101" => n11 <= "0001110110000011";
        when "0110110110" => n11 <= "0001110010000011";
        when "0110110111" => n11 <= "0001110010000011";
        when "0110111000" => n11 <= "0001110010000011";
        when "0110111001" => n11 <= "0001101110000011";
        when "0110111010" => n11 <= "0001101110000010";
        when "0110111011" => n11 <= "0001101010000010";
        when "0110111100" => n11 <= "0001101010000010";
        when "0110111101" => n11 <= "0001101010000010";
        when "0110111110" => n11 <= "0001100110000010";
        when "0110111111" => n11 <= "0001100110000010";
        when "0111000000" => n11 <= "0001100010000010";
        when "0111000001" => n11 <= "0001100010000010";
        when "0111000010" => n11 <= "0001100010000010";
        when "0111000011" => n11 <= "0001011110000010";
        when "0111000100" => n11 <= "0001011110000010";
        when "0111000101" => n11 <= "0001011110000010";
        when "0111000110" => n11 <= "0001011010000010";
        when "0111000111" => n11 <= "0001011010000001";
        when "0111001000" => n11 <= "0001010110000001";
        when "0111001001" => n11 <= "0001010110000001";
        when "0111001010" => n11 <= "0001010110000001";
        when "0111001011" => n11 <= "0001010010000001";
        when "0111001100" => n11 <= "0001010010000001";
        when "0111001101" => n11 <= "0001001110000001";
        when "0111001110" => n11 <= "0001001110000001";
        when "0111001111" => n11 <= "0001001110000001";
        when "0111010000" => n11 <= "0001001010000001";
        when "0111010001" => n11 <= "0001001010000001";
        when "0111010010" => n11 <= "0001001010000001";
        when "0111010011" => n11 <= "0001000110000001";
        when "0111010100" => n11 <= "0001000110000001";
        when "0111010101" => n11 <= "0001000010000001";
        when "0111010110" => n11 <= "0001000010000001";
        when "0111010111" => n11 <= "0001000010000001";
        when "0111011000" => n11 <= "0000111110000000";
        when "0111011001" => n11 <= "0000111110000000";
        when "0111011010" => n11 <= "0000111010000000";
        when "0111011011" => n11 <= "0000111010000000";
        when "0111011100" => n11 <= "0000111010000000";
        when "0111011101" => n11 <= "0000110110000000";
        when "0111011110" => n11 <= "0000110110000000";
        when "0111011111" => n11 <= "0000110010000000";
        when "0111100000" => n11 <= "0000110010000000";
        when "0111100001" => n11 <= "0000110010000000";
        when "0111100010" => n11 <= "0000101110000000";
        when "0111100011" => n11 <= "0000101110000000";
        when "0111100100" => n11 <= "0000101010000000";
        when "0111100101" => n11 <= "0000101010000000";
        when "0111100110" => n11 <= "0000101010000000";
        when "0111100111" => n11 <= "0000100110000000";
        when "0111101000" => n11 <= "0000100110000000";
        when "0111101001" => n11 <= "0000100110000000";
        when "0111101010" => n11 <= "0000100010000000";
        when "0111101011" => n11 <= "0000100010000000";
        when "0111101100" => n11 <= "0000011110000000";
        when "0111101101" => n11 <= "0000011110000000";
        when "0111101110" => n11 <= "0000011110000000";
        when "0111101111" => n11 <= "0000011010000000";
        when "0111110000" => n11 <= "0000011010000000";
        when "0111110001" => n11 <= "0000010110000000";
        when "0111110010" => n11 <= "0000010110000000";
        when "0111110011" => n11 <= "0000010110000000";
        when "0111110100" => n11 <= "0000010010000000";
        when "0111110101" => n11 <= "0000010010000000";
        when "0111110110" => n11 <= "0000001110000000";
        when "0111110111" => n11 <= "0000001110000000";
        when "0111111000" => n11 <= "0000001110000000";
        when "0111111001" => n11 <= "0000001010000000";
        when "0111111010" => n11 <= "0000001010000000";
        when "0111111011" => n11 <= "0000000110000000";
        when "0111111100" => n11 <= "0000000110000000";
        when "0111111101" => n11 <= "0000000110000000";
        when "0111111110" => n11 <= "0000000010000000";
        when "0111111111" => n11 <= "0000000010000000";
        when "1000000000" => n11 <= "0000000010000000";
        when "1000000001" => n11 <= "1111111110000000";
        when "1000000010" => n11 <= "1111111110000000";
        when "1000000011" => n11 <= "1111111010000000";
        when "1000000100" => n11 <= "1111111010000000";
        when "1000000101" => n11 <= "1111111010000000";
        when "1000000110" => n11 <= "1111110110000000";
        when "1000000111" => n11 <= "1111110110000000";
        when "1000001000" => n11 <= "1111110010000000";
        when "1000001001" => n11 <= "1111110010000000";
        when "1000001010" => n11 <= "1111110010000000";
        when "1000001011" => n11 <= "1111101110000000";
        when "1000001100" => n11 <= "1111101110000000";
        when "1000001101" => n11 <= "1111101010000000";
        when "1000001110" => n11 <= "1111101010000000";
        when "1000001111" => n11 <= "1111101010000000";
        when "1000010000" => n11 <= "1111100110000000";
        when "1000010001" => n11 <= "1111100110000000";
        when "1000010010" => n11 <= "1111100010000000";
        when "1000010011" => n11 <= "1111100010000000";
        when "1000010100" => n11 <= "1111100010000000";
        when "1000010101" => n11 <= "1111011110000000";
        when "1000010110" => n11 <= "1111011110000000";
        when "1000010111" => n11 <= "1111011010000000";
        when "1000011000" => n11 <= "1111011010000000";
        when "1000011001" => n11 <= "1111011010000000";
        when "1000011010" => n11 <= "1111010110000000";
        when "1000011011" => n11 <= "1111010110000000";
        when "1000011100" => n11 <= "1111010110000000";
        when "1000011101" => n11 <= "1111010010000000";
        when "1000011110" => n11 <= "1111010010000000";
        when "1000011111" => n11 <= "1111001110000000";
        when "1000100000" => n11 <= "1111001110000000";
        when "1000100001" => n11 <= "1111001110000000";
        when "1000100010" => n11 <= "1111001010000000";
        when "1000100011" => n11 <= "1111001010000000";
        when "1000100100" => n11 <= "1111000110000000";
        when "1000100101" => n11 <= "1111000110000000";
        when "1000100110" => n11 <= "1111000110000000";
        when "1000100111" => n11 <= "1111000010000000";
        when "1000101000" => n11 <= "1111000010000000";
        when "1000101001" => n11 <= "1110111110000001";
        when "1000101010" => n11 <= "1110111110000001";
        when "1000101011" => n11 <= "1110111110000001";
        when "1000101100" => n11 <= "1110111010000001";
        when "1000101101" => n11 <= "1110111010000001";
        when "1000101110" => n11 <= "1110110110000001";
        when "1000101111" => n11 <= "1110110110000001";
        when "1000110000" => n11 <= "1110110110000001";
        when "1000110001" => n11 <= "1110110010000001";
        when "1000110010" => n11 <= "1110110010000001";
        when "1000110011" => n11 <= "1110110010000001";
        when "1000110100" => n11 <= "1110101110000001";
        when "1000110101" => n11 <= "1110101110000001";
        when "1000110110" => n11 <= "1110101010000001";
        when "1000110111" => n11 <= "1110101010000001";
        when "1000111000" => n11 <= "1110101010000001";
        when "1000111001" => n11 <= "1110100110000001";
        when "1000111010" => n11 <= "1110100110000010";
        when "1000111011" => n11 <= "1110100010000010";
        when "1000111100" => n11 <= "1110100010000010";
        when "1000111101" => n11 <= "1110100010000010";
        when "1000111110" => n11 <= "1110011110000010";
        when "1000111111" => n11 <= "1110011110000010";
        when "1001000000" => n11 <= "1110011110000010";
        when "1001000001" => n11 <= "1110011010000010";
        when "1001000010" => n11 <= "1110011010000010";
        when "1001000011" => n11 <= "1110010110000010";
        when "1001000100" => n11 <= "1110010110000010";
        when "1001000101" => n11 <= "1110010110000010";
        when "1001000110" => n11 <= "1110010010000010";
        when "1001000111" => n11 <= "1110010010000011";
        when "1001001000" => n11 <= "1110001110000011";
        when "1001001001" => n11 <= "1110001110000011";
        when "1001001010" => n11 <= "1110001110000011";
        when "1001001011" => n11 <= "1110001010000011";
        when "1001001100" => n11 <= "1110001010000011";
        when "1001001101" => n11 <= "1110001010000011";
        when "1001001110" => n11 <= "1110000110000011";
        when "1001001111" => n11 <= "1110000110000011";
        when "1001010000" => n11 <= "1110000010000011";
        when "1001010001" => n11 <= "1110000010000011";
        when "1001010010" => n11 <= "1110000010000100";
        when "1001010011" => n11 <= "1101111110000100";
        when "1001010100" => n11 <= "1101111110000100";
        when "1001010101" => n11 <= "1101111010000100";
        when "1001010110" => n11 <= "1101111010000100";
        when "1001010111" => n11 <= "1101111010000100";
        when "1001011000" => n11 <= "1101110110000100";
        when "1001011001" => n11 <= "1101110110000100";
        when "1001011010" => n11 <= "1101110110000100";
        when "1001011011" => n11 <= "1101110010000100";
        when "1001011100" => n11 <= "1101110010000101";
        when "1001011101" => n11 <= "1101101110000101";
        when "1001011110" => n11 <= "1101101110000101";
        when "1001011111" => n11 <= "1101101110000101";
        when "1001100000" => n11 <= "1101101010000101";
        when "1001100001" => n11 <= "1101101010000101";
        when "1001100010" => n11 <= "1101101010000101";
        when "1001100011" => n11 <= "1101100110000101";
        when "1001100100" => n11 <= "1101100110000101";
        when "1001100101" => n11 <= "1101100010000110";
        when "1001100110" => n11 <= "1101100010000110";
        when "1001100111" => n11 <= "1101100010000110";
        when "1001101000" => n11 <= "1101011110000110";
        when "1001101001" => n11 <= "1101011110000110";
        when "1001101010" => n11 <= "1101011110000110";
        when "1001101011" => n11 <= "1101011010000110";
        when "1001101100" => n11 <= "1101011010000110";
        when "1001101101" => n11 <= "1101010110000111";
        when "1001101110" => n11 <= "1101010110000111";
        when "1001101111" => n11 <= "1101010110000111";
        when "1001110000" => n11 <= "1101010010000111";
        when "1001110001" => n11 <= "1101010010000111";
        when "1001110010" => n11 <= "1101010010000111";
        when "1001110011" => n11 <= "1101001110000111";
        when "1001110100" => n11 <= "1101001110001000";
        when "1001110101" => n11 <= "1101001110001000";
        when "1001110110" => n11 <= "1101001010001000";
        when "1001110111" => n11 <= "1101001010001000";
        when "1001111000" => n11 <= "1101000110001000";
        when "1001111001" => n11 <= "1101000110001000";
        when "1001111010" => n11 <= "1101000110001000";
        when "1001111011" => n11 <= "1101000010001001";
        when "1001111100" => n11 <= "1101000010001001";
        when "1001111101" => n11 <= "1101000010001001";
        when "1001111110" => n11 <= "1100111110001001";
        when "1001111111" => n11 <= "1100111110001001";
        when "1010000000" => n11 <= "1100111110001001";
        when "1010000001" => n11 <= "1100111010001001";
        when "1010000010" => n11 <= "1100111010001010";
        when "1010000011" => n11 <= "1100110110001010";
        when "1010000100" => n11 <= "1100110110001010";
        when "1010000101" => n11 <= "1100110110001010";
        when "1010000110" => n11 <= "1100110010001010";
        when "1010000111" => n11 <= "1100110010001010";
        when "1010001000" => n11 <= "1100110010001010";
        when "1010001001" => n11 <= "1100101110001011";
        when "1010001010" => n11 <= "1100101110001011";
        when "1010001011" => n11 <= "1100101110001011";
        when "1010001100" => n11 <= "1100101010001011";
        when "1010001101" => n11 <= "1100101010001011";
        when "1010001110" => n11 <= "1100100110001011";
        when "1010001111" => n11 <= "1100100110001100";
        when "1010010000" => n11 <= "1100100110001100";
        when "1010010001" => n11 <= "1100100010001100";
        when "1010010010" => n11 <= "1100100010001100";
        when "1010010011" => n11 <= "1100100010001100";
        when "1010010100" => n11 <= "1100011110001100";
        when "1010010101" => n11 <= "1100011110001101";
        when "1010010110" => n11 <= "1100011110001101";
        when "1010010111" => n11 <= "1100011010001101";
        when "1010011000" => n11 <= "1100011010001101";
        when "1010011001" => n11 <= "1100011010001101";
        when "1010011010" => n11 <= "1100010110001110";
        when "1010011011" => n11 <= "1100010110001110";
        when "1010011100" => n11 <= "1100010110001110";
        when "1010011101" => n11 <= "1100010010001110";
        when "1010011110" => n11 <= "1100010010001110";
        when "1010011111" => n11 <= "1100010010001110";
        when "1010100000" => n11 <= "1100001110001111";
        when "1010100001" => n11 <= "1100001110001111";
        when "1010100010" => n11 <= "1100001010001111";
        when "1010100011" => n11 <= "1100001010001111";
        when "1010100100" => n11 <= "1100001010001111";
        when "1010100101" => n11 <= "1100000110010000";
        when "1010100110" => n11 <= "1100000110010000";
        when "1010100111" => n11 <= "1100000110010000";
        when "1010101000" => n11 <= "1100000010010000";
        when "1010101001" => n11 <= "1100000010010000";
        when "1010101010" => n11 <= "1100000010010001";
        when "1010101011" => n11 <= "1011111110010001";
        when "1010101100" => n11 <= "1011111110010001";
        when "1010101101" => n11 <= "1011111110010001";
        when "1010101110" => n11 <= "1011111010010001";
        when "1010101111" => n11 <= "1011111010010010";
        when "1010110000" => n11 <= "1011111010010010";
        when "1010110001" => n11 <= "1011110110010010";
        when "1010110010" => n11 <= "1011110110010010";
        when "1010110011" => n11 <= "1011110110010010";
        when "1010110100" => n11 <= "1011110010010011";
        when "1010110101" => n11 <= "1011110010010011";
        when "1010110110" => n11 <= "1011110010010011";
        when "1010110111" => n11 <= "1011101110010011";
        when "1010111000" => n11 <= "1011101110010011";
        when "1010111001" => n11 <= "1011101110010100";
        when "1010111010" => n11 <= "1011101010010100";
        when "1010111011" => n11 <= "1011101010010100";
        when "1010111100" => n11 <= "1011101010010100";
        when "1010111101" => n11 <= "1011100110010100";
        when "1010111110" => n11 <= "1011100110010101";
        when "1010111111" => n11 <= "1011100110010101";
        when "1011000000" => n11 <= "1011100010010101";
        when "1011000001" => n11 <= "1011100010010101";
        when "1011000010" => n11 <= "1011100010010110";
        when "1011000011" => n11 <= "1011011110010110";
        when "1011000100" => n11 <= "1011011110010110";
        when "1011000101" => n11 <= "1011011110010110";
        when "1011000110" => n11 <= "1011011010010110";
        when "1011000111" => n11 <= "1011011010010111";
        when "1011001000" => n11 <= "1011011010010111";
        when "1011001001" => n11 <= "1011010110010111";
        when "1011001010" => n11 <= "1011010110010111";
        when "1011001011" => n11 <= "1011010110011000";
        when "1011001100" => n11 <= "1011010110011000";
        when "1011001101" => n11 <= "1011010010011000";
        when "1011001110" => n11 <= "1011010010011000";
        when "1011001111" => n11 <= "1011010010011000";
        when "1011010000" => n11 <= "1011001110011001";
        when "1011010001" => n11 <= "1011001110011001";
        when "1011010010" => n11 <= "1011001110011001";
        when "1011010011" => n11 <= "1011001010011001";
        when "1011010100" => n11 <= "1011001010011010";
        when "1011010101" => n11 <= "1011001010011010";
        when "1011010110" => n11 <= "1011000110011010";
        when "1011010111" => n11 <= "1011000110011010";
        when "1011011000" => n11 <= "1011000110011011";
        when "1011011001" => n11 <= "1011000010011011";
        when "1011011010" => n11 <= "1011000010011011";
        when "1011011011" => n11 <= "1011000010011011";
        when "1011011100" => n11 <= "1011000010011100";
        when "1011011101" => n11 <= "1010111110011100";
        when "1011011110" => n11 <= "1010111110011100";
        when "1011011111" => n11 <= "1010111110011100";
        when "1011100000" => n11 <= "1010111010011101";
        when "1011100001" => n11 <= "1010111010011101";
        when "1011100010" => n11 <= "1010111010011101";
        when "1011100011" => n11 <= "1010110110011101";
        when "1011100100" => n11 <= "1010110110011110";
        when "1011100101" => n11 <= "1010110110011110";
        when "1011100110" => n11 <= "1010110010011110";
        when "1011100111" => n11 <= "1010110010011110";
        when "1011101000" => n11 <= "1010110010011111";
        when "1011101001" => n11 <= "1010110010011111";
        when "1011101010" => n11 <= "1010101110011111";
        when "1011101011" => n11 <= "1010101110011111";
        when "1011101100" => n11 <= "1010101110100000";
        when "1011101101" => n11 <= "1010101010100000";
        when "1011101110" => n11 <= "1010101010100000";
        when "1011101111" => n11 <= "1010101010100000";
        when "1011110000" => n11 <= "1010101010100001";
        when "1011110001" => n11 <= "1010100110100001";
        when "1011110010" => n11 <= "1010100110100001";
        when "1011110011" => n11 <= "1010100110100001";
        when "1011110100" => n11 <= "1010100010100010";
        when "1011110101" => n11 <= "1010100010100010";
        when "1011110110" => n11 <= "1010100010100010";
        when "1011110111" => n11 <= "1010100010100011";
        when "1011111000" => n11 <= "1010011110100011";
        when "1011111001" => n11 <= "1010011110100011";
        when "1011111010" => n11 <= "1010011110100011";
        when "1011111011" => n11 <= "1010011010100100";
        when "1011111100" => n11 <= "1010011010100100";
        when "1011111101" => n11 <= "1010011010100100";
        when "1011111110" => n11 <= "1010011010100100";
        when "1011111111" => n11 <= "1010010110100101";
        when "1100000000" => n11 <= "1010010110100101";
        when "1100000001" => n11 <= "1010010110100101";
        when "1100000010" => n11 <= "1010010010100110";
        when "1100000011" => n11 <= "1010010010100110";
        when "1100000100" => n11 <= "1010010010100110";
        when "1100000101" => n11 <= "1010010010100110";
        when "1100000110" => n11 <= "1010001110100111";
        when "1100000111" => n11 <= "1010001110100111";
        when "1100001000" => n11 <= "1010001110100111";
        when "1100001001" => n11 <= "1010001110101000";
        when "1100001010" => n11 <= "1010001010101000";
        when "1100001011" => n11 <= "1010001010101000";
        when "1100001100" => n11 <= "1010001010101000";
        when "1100001101" => n11 <= "1010000110101001";
        when "1100001110" => n11 <= "1010000110101001";
        when "1100001111" => n11 <= "1010000110101001";
        when "1100010000" => n11 <= "1010000110101010";
        when "1100010001" => n11 <= "1010000010101010";
        when "1100010010" => n11 <= "1010000010101010";
        when "1100010011" => n11 <= "1010000010101010";
        when "1100010100" => n11 <= "1010000010101011";
        when "1100010101" => n11 <= "1001111110101011";
        when "1100010110" => n11 <= "1001111110101011";
        when "1100010111" => n11 <= "1001111110101100";
        when "1100011000" => n11 <= "1001111110101100";
        when "1100011001" => n11 <= "1001111010101100";
        when "1100011010" => n11 <= "1001111010101100";
        when "1100011011" => n11 <= "1001111010101101";
        when "1100011100" => n11 <= "1001111010101101";
        when "1100011101" => n11 <= "1001110110101101";
        when "1100011110" => n11 <= "1001110110101110";
        when "1100011111" => n11 <= "1001110110101110";
        when "1100100000" => n11 <= "1001110110101110";
        when "1100100001" => n11 <= "1001110010101111";
        when "1100100010" => n11 <= "1001110010101111";
        when "1100100011" => n11 <= "1001110010101111";
        when "1100100100" => n11 <= "1001110010110000";
        when "1100100101" => n11 <= "1001101110110000";
        when "1100100110" => n11 <= "1001101110110000";
        when "1100100111" => n11 <= "1001101110110000";
        when "1100101000" => n11 <= "1001101110110001";
        when "1100101001" => n11 <= "1001101010110001";
        when "1100101010" => n11 <= "1001101010110001";
        when "1100101011" => n11 <= "1001101010110010";
        when "1100101100" => n11 <= "1001101010110010";
        when "1100101101" => n11 <= "1001100110110010";
        when "1100101110" => n11 <= "1001100110110011";
        when "1100101111" => n11 <= "1001100110110011";
        when "1100110000" => n11 <= "1001100110110011";
        when "1100110001" => n11 <= "1001100010110100";
        when "1100110010" => n11 <= "1001100010110100";
        when "1100110011" => n11 <= "1001100010110100";
        when "1100110100" => n11 <= "1001100010110101";
        when "1100110101" => n11 <= "1001100010110101";
        when "1100110110" => n11 <= "1001011110110101";
        when "1100110111" => n11 <= "1001011110110101";
        when "1100111000" => n11 <= "1001011110110110";
        when "1100111001" => n11 <= "1001011110110110";
        when "1100111010" => n11 <= "1001011010110110";
        when "1100111011" => n11 <= "1001011010110111";
        when "1100111100" => n11 <= "1001011010110111";
        when "1100111101" => n11 <= "1001011010110111";
        when "1100111110" => n11 <= "1001011010111000";
        when "1100111111" => n11 <= "1001010110111000";
        when "1101000000" => n11 <= "1001010110111000";
        when "1101000001" => n11 <= "1001010110111001";
        when "1101000010" => n11 <= "1001010110111001";
        when "1101000011" => n11 <= "1001010010111001";
        when "1101000100" => n11 <= "1001010010111010";
        when "1101000101" => n11 <= "1001010010111010";
        when "1101000110" => n11 <= "1001010010111010";
        when "1101000111" => n11 <= "1001010010111011";
        when "1101001000" => n11 <= "1001001110111011";
        when "1101001001" => n11 <= "1001001110111011";
        when "1101001010" => n11 <= "1001001110111100";
        when "1101001011" => n11 <= "1001001110111100";
        when "1101001100" => n11 <= "1001001110111100";
        when "1101001101" => n11 <= "1001001010111101";
        when "1101001110" => n11 <= "1001001010111101";
        when "1101001111" => n11 <= "1001001010111101";
        when "1101010000" => n11 <= "1001001010111110";
        when "1101010001" => n11 <= "1001001010111110";
        when "1101010010" => n11 <= "1001000110111110";
        when "1101010011" => n11 <= "1001000110111111";
        when "1101010100" => n11 <= "1001000110111111";
        when "1101010101" => n11 <= "1001000110111111";
        when "1101010110" => n11 <= "1001000111000000";
        when "1101010111" => n11 <= "1001000011000000";
        when "1101011000" => n11 <= "1001000011000000";
        when "1101011001" => n11 <= "1001000011000001";
        when "1101011010" => n11 <= "1001000011000001";
        when "1101011011" => n11 <= "1001000011000001";
        when "1101011100" => n11 <= "1000111111000010";
        when "1101011101" => n11 <= "1000111111000010";
        when "1101011110" => n11 <= "1000111111000010";
        when "1101011111" => n11 <= "1000111111000011";
        when "1101100000" => n11 <= "1000111111000011";
        when "1101100001" => n11 <= "1000111011000100";
        when "1101100010" => n11 <= "1000111011000100";
        when "1101100011" => n11 <= "1000111011000100";
        when "1101100100" => n11 <= "1000111011000101";
        when "1101100101" => n11 <= "1000111011000101";
        when "1101100110" => n11 <= "1000111011000101";
        when "1101100111" => n11 <= "1000110111000110";
        when "1101101000" => n11 <= "1000110111000110";
        when "1101101001" => n11 <= "1000110111000110";
        when "1101101010" => n11 <= "1000110111000111";
        when "1101101011" => n11 <= "1000110111000111";
        when "1101101100" => n11 <= "1000110011000111";
        when "1101101101" => n11 <= "1000110011001000";
        when "1101101110" => n11 <= "1000110011001000";
        when "1101101111" => n11 <= "1000110011001000";
        when "1101110000" => n11 <= "1000110011001001";
        when "1101110001" => n11 <= "1000110011001001";
        when "1101110010" => n11 <= "1000101111001001";
        when "1101110011" => n11 <= "1000101111001010";
        when "1101110100" => n11 <= "1000101111001010";
        when "1101110101" => n11 <= "1000101111001011";
        when "1101110110" => n11 <= "1000101111001011";
        when "1101110111" => n11 <= "1000101111001011";
        when "1101111000" => n11 <= "1000101011001100";
        when "1101111001" => n11 <= "1000101011001100";
        when "1101111010" => n11 <= "1000101011001100";
        when "1101111011" => n11 <= "1000101011001101";
        when "1101111100" => n11 <= "1000101011001101";
        when "1101111101" => n11 <= "1000101011001101";
        when "1101111110" => n11 <= "1000101011001110";
        when "1101111111" => n11 <= "1000100111001110";
        when "1110000000" => n11 <= "1000100111001111";
        when "1110000001" => n11 <= "1000100111001111";
        when "1110000010" => n11 <= "1000100111001111";
        when "1110000011" => n11 <= "1000100111010000";
        when "1110000100" => n11 <= "1000100111010000";
        when "1110000101" => n11 <= "1000100111010000";
        when "1110000110" => n11 <= "1000100011010001";
        when "1110000111" => n11 <= "1000100011010001";
        when "1110001000" => n11 <= "1000100011010001";
        when "1110001001" => n11 <= "1000100011010010";
        when "1110001010" => n11 <= "1000100011010010";
        when "1110001011" => n11 <= "1000100011010011";
        when "1110001100" => n11 <= "1000100011010011";
        when "1110001101" => n11 <= "1000011111010011";
        when "1110001110" => n11 <= "1000011111010100";
        when "1110001111" => n11 <= "1000011111010100";
        when "1110010000" => n11 <= "1000011111010100";
        when "1110010001" => n11 <= "1000011111010101";
        when "1110010010" => n11 <= "1000011111010101";
        when "1110010011" => n11 <= "1000011111010101";
        when "1110010100" => n11 <= "1000011011010110";
        when "1110010101" => n11 <= "1000011011010110";
        when "1110010110" => n11 <= "1000011011010111";
        when "1110010111" => n11 <= "1000011011010111";
        when "1110011000" => n11 <= "1000011011010111";
        when "1110011001" => n11 <= "1000011011011000";
        when "1110011010" => n11 <= "1000011011011000";
        when "1110011011" => n11 <= "1000011011011000";
        when "1110011100" => n11 <= "1000010111011001";
        when "1110011101" => n11 <= "1000010111011001";
        when "1110011110" => n11 <= "1000010111011010";
        when "1110011111" => n11 <= "1000010111011010";
        when "1110100000" => n11 <= "1000010111011010";
        when "1110100001" => n11 <= "1000010111011011";
        when "1110100010" => n11 <= "1000010111011011";
        when "1110100011" => n11 <= "1000010111011011";
        when "1110100100" => n11 <= "1000010111011100";
        when "1110100101" => n11 <= "1000010011011100";
        when "1110100110" => n11 <= "1000010011011101";
        when "1110100111" => n11 <= "1000010011011101";
        when "1110101000" => n11 <= "1000010011011101";
        when "1110101001" => n11 <= "1000010011011110";
        when "1110101010" => n11 <= "1000010011011110";
        when "1110101011" => n11 <= "1000010011011110";
        when "1110101100" => n11 <= "1000010011011111";
        when "1110101101" => n11 <= "1000010011011111";
        when "1110101110" => n11 <= "1000010011100000";
        when "1110101111" => n11 <= "1000001111100000";
        when "1110110000" => n11 <= "1000001111100000";
        when "1110110001" => n11 <= "1000001111100001";
        when "1110110010" => n11 <= "1000001111100001";
        when "1110110011" => n11 <= "1000001111100010";
        when "1110110100" => n11 <= "1000001111100010";
        when "1110110101" => n11 <= "1000001111100010";
        when "1110110110" => n11 <= "1000001111100011";
        when "1110110111" => n11 <= "1000001111100011";
        when "1110111000" => n11 <= "1000001111100011";
        when "1110111001" => n11 <= "1000001111100100";
        when "1110111010" => n11 <= "1000001011100100";
        when "1110111011" => n11 <= "1000001011100101";
        when "1110111100" => n11 <= "1000001011100101";
        when "1110111101" => n11 <= "1000001011100101";
        when "1110111110" => n11 <= "1000001011100110";
        when "1110111111" => n11 <= "1000001011100110";
        when "1111000000" => n11 <= "1000001011100111";
        when "1111000001" => n11 <= "1000001011100111";
        when "1111000010" => n11 <= "1000001011100111";
        when "1111000011" => n11 <= "1000001011101000";
        when "1111000100" => n11 <= "1000001011101000";
        when "1111000101" => n11 <= "1000001011101000";
        when "1111000110" => n11 <= "1000001011101001";
        when "1111000111" => n11 <= "1000000111101001";
        when "1111001000" => n11 <= "1000000111101010";
        when "1111001001" => n11 <= "1000000111101010";
        when "1111001010" => n11 <= "1000000111101010";
        when "1111001011" => n11 <= "1000000111101011";
        when "1111001100" => n11 <= "1000000111101011";
        when "1111001101" => n11 <= "1000000111101100";
        when "1111001110" => n11 <= "1000000111101100";
        when "1111001111" => n11 <= "1000000111101100";
        when "1111010000" => n11 <= "1000000111101101";
        when "1111010001" => n11 <= "1000000111101101";
        when "1111010010" => n11 <= "1000000111101101";
        when "1111010011" => n11 <= "1000000111101110";
        when "1111010100" => n11 <= "1000000111101110";
        when "1111010101" => n11 <= "1000000111101111";
        when "1111010110" => n11 <= "1000000111101111";
        when "1111010111" => n11 <= "1000000111101111";
        when "1111011000" => n11 <= "1000000011110000";
        when "1111011001" => n11 <= "1000000011110000";
        when "1111011010" => n11 <= "1000000011110001";
        when "1111011011" => n11 <= "1000000011110001";
        when "1111011100" => n11 <= "1000000011110001";
        when "1111011101" => n11 <= "1000000011110010";
        when "1111011110" => n11 <= "1000000011110010";
        when "1111011111" => n11 <= "1000000011110011";
        when "1111100000" => n11 <= "1000000011110011";
        when "1111100001" => n11 <= "1000000011110011";
        when "1111100010" => n11 <= "1000000011110100";
        when "1111100011" => n11 <= "1000000011110100";
        when "1111100100" => n11 <= "1000000011110101";
        when "1111100101" => n11 <= "1000000011110101";
        when "1111100110" => n11 <= "1000000011110101";
        when "1111100111" => n11 <= "1000000011110110";
        when "1111101000" => n11 <= "1000000011110110";
        when "1111101001" => n11 <= "1000000011110110";
        when "1111101010" => n11 <= "1000000011110111";
        when "1111101011" => n11 <= "1000000011110111";
        when "1111101100" => n11 <= "1000000011111000";
        when "1111101101" => n11 <= "1000000011111000";
        when "1111101110" => n11 <= "1000000011111000";
        when "1111101111" => n11 <= "1000000011111001";
        when "1111110000" => n11 <= "1000000011111001";
        when "1111110001" => n11 <= "1000000011111010";
        when "1111110010" => n11 <= "1000000011111010";
        when "1111110011" => n11 <= "1000000011111010";
        when "1111110100" => n11 <= "1000000011111011";
        when "1111110101" => n11 <= "1000000011111011";
        when "1111110110" => n11 <= "1000000011111100";
        when "1111110111" => n11 <= "1000000011111100";
        when "1111111000" => n11 <= "1000000011111100";
        when "1111111001" => n11 <= "1000000011111101";
        when "1111111010" => n11 <= "1000000011111101";
        when "1111111011" => n11 <= "1000000011111110";
        when "1111111100" => n11 <= "1000000011111110";
        when "1111111101" => n11 <= "1000000011111110";
        when "1111111110" => n11 <= "1000000011111111";
        when "1111111111" => n11 <= "1000000011111111";
        when others => n11 <= "XXXXXXXXXXXXXXXX";
      end case;
    end if;
  end if;
end process;
n12 <= n11(15 downto 15) &
  n11(14 downto 14) &
  n11(13 downto 13) &
  n11(12 downto 12) &
  n11(11 downto 11) &
  n11(10 downto 10) &
  n11(9 downto 9) &
  n11(8 downto 8);
n13 <= n11(7 downto 7) &
  n11(6 downto 6) &
  n11(5 downto 5) &
  n11(4 downto 4) &
  n11(3 downto 3) &
  n11(2 downto 2) &
  n11(1 downto 1) &
  n11(0 downto 0);
n14 <= unsigned(signed(n5) * signed(n12));
n15 <= n14(14 downto 14) &
  n14(13 downto 13) &
  n14(12 downto 12) &
  n14(11 downto 11) &
  n14(10 downto 10) &
  n14(9 downto 9) &
  n14(8 downto 8) &
  n14(7 downto 7);
process (clock_c) begin
  if rising_edge(clock_c) then
    if i5 = "1" then
      n16 <= "00000000";
    elsif i4 = "1" then
      n16 <= n15;
    end if;
  end if;
end process;
n17 <= unsigned(signed(n6) * signed(n13));
n18 <= n17(14 downto 14) &
  n17(13 downto 13) &
  n17(12 downto 12) &
  n17(11 downto 11) &
  n17(10 downto 10) &
  n17(9 downto 9) &
  n17(8 downto 8) &
  n17(7 downto 7);
process (clock_c) begin
  if rising_edge(clock_c) then
    if i5 = "1" then
      n19 <= "00000000";
    elsif i4 = "1" then
      n19 <= n18;
    end if;
  end if;
end process;
n20 <= n16 - n19;
process (clock_c) begin
  if rising_edge(clock_c) then
    if i5 = "1" then
      n21 <= "00000000";
    elsif i4 = "1" then
      n21 <= n20;
    end if;
  end if;
end process;
n22 <= unsigned(signed(n5) * signed(n13));
n23 <= n22(14 downto 14) &
  n22(13 downto 13) &
  n22(12 downto 12) &
  n22(11 downto 11) &
  n22(10 downto 10) &
  n22(9 downto 9) &
  n22(8 downto 8) &
  n22(7 downto 7);
process (clock_c) begin
  if rising_edge(clock_c) then
    if i5 = "1" then
      n24 <= "00000000";
    elsif i4 = "1" then
      n24 <= n23;
    end if;
  end if;
end process;
n25 <= unsigned(signed(n6) * signed(n12));
n26 <= n25(14 downto 14) &
  n25(13 downto 13) &
  n25(12 downto 12) &
  n25(11 downto 11) &
  n25(10 downto 10) &
  n25(9 downto 9) &
  n25(8 downto 8) &
  n25(7 downto 7);
process (clock_c) begin
  if rising_edge(clock_c) then
    if i5 = "1" then
      n27 <= "00000000";
    elsif i4 = "1" then
      n27 <= n26;
    end if;
  end if;
end process;
n28 <= n24 + n27;
process (clock_c) begin
  if rising_edge(clock_c) then
    if i5 = "1" then
      n29 <= "00000000";
    elsif i4 = "1" then
      n29 <= n28;
    end if;
  end if;
end process;
n30 <= n8 + n21;
n31 <= n10 + n29;
n32 <= n30 & n31;
process (clock_c) begin
  if rising_edge(clock_c) then
    if i5 = "1" then
      n33 <= "0000000000000000";
    elsif i4 = "1" then
      n33 <= n32;
    end if;
  end if;
end process;
n34 <= n8 - n21;
n35 <= n10 - n29;
n36 <= n34 & n35;
process (clock_c) begin
  if rising_edge(clock_c) then
    if i5 = "1" then
      n37 <= "0000000000000000";
    elsif i4 = "1" then
      n37 <= n36;
    end if;
  end if;
end process;
o2 <= n37;
o1 <= n33;
end architecture rtl;

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
entity cf_fft_2048_8_23 is
port (
clock_c : in std_logic;
i1 : in  unsigned(0 downto 0);
i2 : in  unsigned(15 downto 0);
i3 : in  unsigned(15 downto 0);
i4 : in  unsigned(0 downto 0);
i5 : in  unsigned(0 downto 0);
o1 : out unsigned(0 downto 0);
o2 : out unsigned(15 downto 0);
o3 : out unsigned(15 downto 0));
end entity cf_fft_2048_8_23;
architecture rtl of cf_fft_2048_8_23 is
signal n1 : unsigned(9 downto 0);
signal n2 : unsigned(31 downto 0);
signal n3 : unsigned(0 downto 0) := "0";
signal n4 : unsigned(0 downto 0) := "0";
signal n5 : unsigned(0 downto 0) := "0";
signal n6 : unsigned(0 downto 0) := "0";
signal n7 : unsigned(8 downto 0);
signal n8 : unsigned(8 downto 0) := "000000000";
signal n9 : unsigned(8 downto 0) := "000000000";
signal n10 : unsigned(8 downto 0) := "000000000";
signal n11 : unsigned(8 downto 0) := "000000000";
signal n12 : unsigned(0 downto 0);
signal n13 : unsigned(0 downto 0) := "0";
signal n14 : unsigned(0 downto 0) := "0";
signal n15 : unsigned(0 downto 0) := "0";
signal n16 : unsigned(0 downto 0) := "0";
signal n17 : unsigned(0 downto 0);
signal n18 : unsigned(1 downto 0);
signal n19 : unsigned(15 downto 0);
signal n20 : unsigned(15 downto 0);
signal n21 : unsigned(15 downto 0);
signal n22 : unsigned(15 downto 0);
signal n23 : unsigned(15 downto 0);
signal n24 : unsigned(15 downto 0);
signal s25_1 : unsigned(15 downto 0);
signal s25_2 : unsigned(15 downto 0);
signal s26_1 : unsigned(0 downto 0);
signal s27_1 : unsigned(31 downto 0);
signal s28_1 : unsigned(0 downto 0);
signal s28_2 : unsigned(0 downto 0);
signal s28_3 : unsigned(31 downto 0);
signal s29_1 : unsigned(9 downto 0);
signal s29_2 : unsigned(0 downto 0);
component cf_fft_2048_8_24 is
port (
clock_c : in std_logic;
i1 : in  unsigned(15 downto 0);
i2 : in  unsigned(15 downto 0);
i3 : in  unsigned(9 downto 0);
i4 : in  unsigned(0 downto 0);
i5 : in  unsigned(0 downto 0);
o1 : out unsigned(15 downto 0);
o2 : out unsigned(15 downto 0));
end component cf_fft_2048_8_24;
component cf_fft_2048_8_35 is
port (
clock_c : in std_logic;
i1 : in  unsigned(1 downto 0);
i2 : in  unsigned(0 downto 0);
i3 : in  unsigned(0 downto 0);
o1 : out unsigned(0 downto 0));
end component cf_fft_2048_8_35;
component cf_fft_2048_8_31 is
port (
clock_c : in std_logic;
i1 : in  unsigned(31 downto 0);
i2 : in  unsigned(0 downto 0);
i3 : in  unsigned(8 downto 0);
i4 : in  unsigned(0 downto 0);
i5 : in  unsigned(0 downto 0);
i6 : in  unsigned(0 downto 0);
o1 : out unsigned(31 downto 0));
end component cf_fft_2048_8_31;
component cf_fft_2048_8_30 is
port (
clock_c : in std_logic;
i1 : in  unsigned(31 downto 0);
i2 : in  unsigned(0 downto 0);
i3 : in  unsigned(8 downto 0);
i4 : in  unsigned(0 downto 0);
i5 : in  unsigned(0 downto 0);
i6 : in  unsigned(0 downto 0);
o1 : out unsigned(0 downto 0);
o2 : out unsigned(0 downto 0);
o3 : out unsigned(31 downto 0));
end component cf_fft_2048_8_30;
component cf_fft_2048_8_26 is
port (
clock_c : in std_logic;
i1 : in  unsigned(0 downto 0);
i2 : in  unsigned(0 downto 0);
i3 : in  unsigned(0 downto 0);
o1 : out unsigned(9 downto 0);
o2 : out unsigned(0 downto 0));
end component cf_fft_2048_8_26;
begin
n1 <= s29_1(9 downto 9) &
  s29_1(8 downto 8) &
  s29_1(7 downto 7) &
  s29_1(6 downto 6) &
  s29_1(5 downto 5) &
  s29_1(4 downto 4) &
  s29_1(3 downto 3) &
  s29_1(2 downto 2) &
  s29_1(1 downto 1) &
  s29_1(0 downto 0);
n2 <= s25_1 & s25_2;
process (clock_c) begin
  if rising_edge(clock_c) then
    if i5 = "1" then
      n3 <= "0";
    elsif i4 = "1" then
      n3 <= s29_2;
    end if;
  end if;
end process;
process (clock_c) begin
  if rising_edge(clock_c) then
    if i5 = "1" then
      n4 <= "0";
    elsif i4 = "1" then
      n4 <= n3;
    end if;
  end if;
end process;
process (clock_c) begin
  if rising_edge(clock_c) then
    if i5 = "1" then
      n5 <= "0";
    elsif i4 = "1" then
      n5 <= n4;
    end if;
  end if;
end process;
process (clock_c) begin
  if rising_edge(clock_c) then
    if i5 = "1" then
      n6 <= "0";
    elsif i4 = "1" then
      n6 <= n5;
    end if;
  end if;
end process;
n7 <= s29_1(9 downto 9) &
  s29_1(8 downto 8) &
  s29_1(7 downto 7) &
  s29_1(6 downto 6) &
  s29_1(5 downto 5) &
  s29_1(4 downto 4) &
  s29_1(3 downto 3) &
  s29_1(2 downto 2) &
  s29_1(1 downto 1);
process (clock_c) begin
  if rising_edge(clock_c) then
    if i5 = "1" then
      n8 <= "000000000";
    elsif i4 = "1" then
      n8 <= n7;
    end if;
  end if;
end process;
process (clock_c) begin
  if rising_edge(clock_c) then
    if i5 = "1" then
      n9 <= "000000000";
    elsif i4 = "1" then
      n9 <= n8;
    end if;
  end if;
end process;
process (clock_c) begin
  if rising_edge(clock_c) then
    if i5 = "1" then
      n10 <= "000000000";
    elsif i4 = "1" then
      n10 <= n9;
    end if;
  end if;
end process;
process (clock_c) begin
  if rising_edge(clock_c) then
    if i5 = "1" then
      n11 <= "000000000";
    elsif i4 = "1" then
      n11 <= n10;
    end if;
  end if;
end process;
n12 <= s29_1(0 downto 0);
process (clock_c) begin
  if rising_edge(clock_c) then
    if i5 = "1" then
      n13 <= "0";
    elsif i4 = "1" then
      n13 <= n12;
    end if;
  end if;
end process;
process (clock_c) begin
  if rising_edge(clock_c) then
    if i5 = "1" then
      n14 <= "0";
    elsif i4 = "1" then
      n14 <= n13;
    end if;
  end if;
end process;
process (clock_c) begin
  if rising_edge(clock_c) then
    if i5 = "1" then
      n15 <= "0";
    elsif i4 = "1" then
      n15 <= n14;
    end if;
  end if;
end process;
process (clock_c) begin
  if rising_edge(clock_c) then
    if i5 = "1" then
      n16 <= "0";
    elsif i4 = "1" then
      n16 <= n15;
    end if;
  end if;
end process;
n17 <= not n16;
n18 <= s28_2 & s28_1;
n19 <= s28_3(31 downto 31) &
  s28_3(30 downto 30) &
  s28_3(29 downto 29) &
  s28_3(28 downto 28) &
  s28_3(27 downto 27) &
  s28_3(26 downto 26) &
  s28_3(25 downto 25) &
  s28_3(24 downto 24) &
  s28_3(23 downto 23) &
  s28_3(22 downto 22) &
  s28_3(21 downto 21) &
  s28_3(20 downto 20) &
  s28_3(19 downto 19) &
  s28_3(18 downto 18) &
  s28_3(17 downto 17) &
  s28_3(16 downto 16);
n20 <= s28_3(15 downto 15) &
  s28_3(14 downto 14) &
  s28_3(13 downto 13) &
  s28_3(12 downto 12) &
  s28_3(11 downto 11) &
  s28_3(10 downto 10) &
  s28_3(9 downto 9) &
  s28_3(8 downto 8) &
  s28_3(7 downto 7) &
  s28_3(6 downto 6) &
  s28_3(5 downto 5) &
  s28_3(4 downto 4) &
  s28_3(3 downto 3) &
  s28_3(2 downto 2) &
  s28_3(1 downto 1) &
  s28_3(0 downto 0);
n21 <= s27_1(31 downto 31) &
  s27_1(30 downto 30) &
  s27_1(29 downto 29) &
  s27_1(28 downto 28) &
  s27_1(27 downto 27) &
  s27_1(26 downto 26) &
  s27_1(25 downto 25) &
  s27_1(24 downto 24) &
  s27_1(23 downto 23) &
  s27_1(22 downto 22) &
  s27_1(21 downto 21) &
  s27_1(20 downto 20) &
  s27_1(19 downto 19) &
  s27_1(18 downto 18) &
  s27_1(17 downto 17) &
  s27_1(16 downto 16);
n22 <= s27_1(15 downto 15) &
  s27_1(14 downto 14) &
  s27_1(13 downto 13) &
  s27_1(12 downto 12) &
  s27_1(11 downto 11) &
  s27_1(10 downto 10) &
  s27_1(9 downto 9) &
  s27_1(8 downto 8) &
  s27_1(7 downto 7) &
  s27_1(6 downto 6) &
  s27_1(5 downto 5) &
  s27_1(4 downto 4) &
  s27_1(3 downto 3) &
  s27_1(2 downto 2) &
  s27_1(1 downto 1) &
  s27_1(0 downto 0);
n23 <= n20 when s26_1 = "1" else n19;
n24 <= n22 when s26_1 = "1" else n21;
s25 : cf_fft_2048_8_24 port map (clock_c, i2, i3, n1, i4, i5, s25_1, s25_2);
s26 : cf_fft_2048_8_35 port map (clock_c, n18, i4, i5, s26_1);
s27 : cf_fft_2048_8_31 port map (clock_c, n2, n6, n11, n16, i4, i5, s27_1);
s28 : cf_fft_2048_8_30 port map (clock_c, n2, n6, n11, n17, i4, i5, s28_1, s28_2, s28_3);
s29 : cf_fft_2048_8_26 port map (clock_c, i1, i4, i5, s29_1, s29_2);
o3 <= n24;
o2 <= n23;
o1 <= s28_1;
end architecture rtl;

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
entity cf_fft_2048_8_22 is
port (
clock_c : in std_logic;
i1 : in  unsigned(15 downto 0);
i2 : in  unsigned(15 downto 0);
i3 : in  unsigned(8 downto 0);
i4 : in  unsigned(0 downto 0);
i5 : in  unsigned(0 downto 0);
o1 : out unsigned(15 downto 0);
o2 : out unsigned(15 downto 0));
end entity cf_fft_2048_8_22;
architecture rtl of cf_fft_2048_8_22 is
signal n1 : unsigned(15 downto 0) := "0000000000000000";
signal n2 : unsigned(7 downto 0);
signal n3 : unsigned(7 downto 0);
signal n4 : unsigned(15 downto 0) := "0000000000000000";
signal n5 : unsigned(7 downto 0);
signal n6 : unsigned(7 downto 0);
signal n7 : unsigned(7 downto 0) := "00000000";
signal n8 : unsigned(7 downto 0) := "00000000";
signal n9 : unsigned(7 downto 0) := "00000000";
signal n10 : unsigned(7 downto 0) := "00000000";
signal n11 : unsigned(15 downto 0) := "0000000000000000";
signal n12 : unsigned(7 downto 0);
signal n13 : unsigned(7 downto 0);
signal n14 : unsigned(15 downto 0);
signal n15 : unsigned(7 downto 0);
signal n16 : unsigned(7 downto 0) := "00000000";
signal n17 : unsigned(15 downto 0);
signal n18 : unsigned(7 downto 0);
signal n19 : unsigned(7 downto 0) := "00000000";
signal n20 : unsigned(7 downto 0);
signal n21 : unsigned(7 downto 0) := "00000000";
signal n22 : unsigned(15 downto 0);
signal n23 : unsigned(7 downto 0);
signal n24 : unsigned(7 downto 0) := "00000000";
signal n25 : unsigned(15 downto 0);
signal n26 : unsigned(7 downto 0);
signal n27 : unsigned(7 downto 0) := "00000000";
signal n28 : unsigned(7 downto 0);
signal n29 : unsigned(7 downto 0) := "00000000";
signal n30 : unsigned(7 downto 0);
signal n31 : unsigned(7 downto 0);
signal n32 : unsigned(15 downto 0);
signal n33 : unsigned(15 downto 0) := "0000000000000000";
signal n34 : unsigned(7 downto 0);
signal n35 : unsigned(7 downto 0);
signal n36 : unsigned(15 downto 0);
signal n37 : unsigned(15 downto 0) := "0000000000000000";
begin
process (clock_c) begin
  if rising_edge(clock_c) then
    if i5 = "1" then
      n1 <= "0000000000000000";
    elsif i4 = "1" then
      n1 <= i1;
    end if;
  end if;
end process;
n2 <= n1(15 downto 15) &
  n1(14 downto 14) &
  n1(13 downto 13) &
  n1(12 downto 12) &
  n1(11 downto 11) &
  n1(10 downto 10) &
  n1(9 downto 9) &
  n1(8 downto 8);
n3 <= n1(7 downto 7) &
  n1(6 downto 6) &
  n1(5 downto 5) &
  n1(4 downto 4) &
  n1(3 downto 3) &
  n1(2 downto 2) &
  n1(1 downto 1) &
  n1(0 downto 0);
process (clock_c) begin
  if rising_edge(clock_c) then
    if i5 = "1" then
      n4 <= "0000000000000000";
    elsif i4 = "1" then
      n4 <= i2;
    end if;
  end if;
end process;
n5 <= n4(15 downto 15) &
  n4(14 downto 14) &
  n4(13 downto 13) &
  n4(12 downto 12) &
  n4(11 downto 11) &
  n4(10 downto 10) &
  n4(9 downto 9) &
  n4(8 downto 8);
n6 <= n4(7 downto 7) &
  n4(6 downto 6) &
  n4(5 downto 5) &
  n4(4 downto 4) &
  n4(3 downto 3) &
  n4(2 downto 2) &
  n4(1 downto 1) &
  n4(0 downto 0);
process (clock_c) begin
  if rising_edge(clock_c) then
    if i5 = "1" then
      n7 <= "00000000";
    elsif i4 = "1" then
      n7 <= n2;
    end if;
  end if;
end process;
process (clock_c) begin
  if rising_edge(clock_c) then
    if i5 = "1" then
      n8 <= "00000000";
    elsif i4 = "1" then
      n8 <= n7;
    end if;
  end if;
end process;
process (clock_c) begin
  if rising_edge(clock_c) then
    if i5 = "1" then
      n9 <= "00000000";
    elsif i4 = "1" then
      n9 <= n3;
    end if;
  end if;
end process;
process (clock_c) begin
  if rising_edge(clock_c) then
    if i5 = "1" then
      n10 <= "00000000";
    elsif i4 = "1" then
      n10 <= n9;
    end if;
  end if;
end process;
process (clock_c) begin
  if rising_edge(clock_c) then 
    if i4 = "1" then
      case i3 is
        when "000000000" => n11 <= "0111111100000000";
        when "000000001" => n11 <= "0111111111111111";
        when "000000010" => n11 <= "0111111111111110";
        when "000000011" => n11 <= "0111111111111101";
        when "000000100" => n11 <= "0111111111111100";
        when "000000101" => n11 <= "0111111111111100";
        when "000000110" => n11 <= "0111111111111011";
        when "000000111" => n11 <= "0111111111111010";
        when "000001000" => n11 <= "0111111111111001";
        when "000001001" => n11 <= "0111111111111000";
        when "000001010" => n11 <= "0111111111111000";
        when "000001011" => n11 <= "0111111111110111";
        when "000001100" => n11 <= "0111111111110110";
        when "000001101" => n11 <= "0111111111110101";
        when "000001110" => n11 <= "0111111111110101";
        when "000001111" => n11 <= "0111111111110100";
        when "000010000" => n11 <= "0111111111110011";
        when "000010001" => n11 <= "0111111111110010";
        when "000010010" => n11 <= "0111111111110001";
        when "000010011" => n11 <= "0111111111110001";
        when "000010100" => n11 <= "0111111111110000";
        when "000010101" => n11 <= "0111111011101111";
        when "000010110" => n11 <= "0111111011101110";
        when "000010111" => n11 <= "0111111011101101";
        when "000011000" => n11 <= "0111111011101101";
        when "000011001" => n11 <= "0111111011101100";
        when "000011010" => n11 <= "0111111011101011";
        when "000011011" => n11 <= "0111111011101010";
        when "000011100" => n11 <= "0111111011101010";
        when "000011101" => n11 <= "0111110111101001";
        when "000011110" => n11 <= "0111110111101000";
        when "000011111" => n11 <= "0111110111100111";
        when "000100000" => n11 <= "0111110111100111";
        when "000100001" => n11 <= "0111110111100110";
        when "000100010" => n11 <= "0111110111100101";
        when "000100011" => n11 <= "0111110111100100";
        when "000100100" => n11 <= "0111110011100011";
        when "000100101" => n11 <= "0111110011100011";
        when "000100110" => n11 <= "0111110011100010";
        when "000100111" => n11 <= "0111110011100001";
        when "000101000" => n11 <= "0111110011100000";
        when "000101001" => n11 <= "0111101111100000";
        when "000101010" => n11 <= "0111101111011111";
        when "000101011" => n11 <= "0111101111011110";
        when "000101100" => n11 <= "0111101111011101";
        when "000101101" => n11 <= "0111101111011101";
        when "000101110" => n11 <= "0111101011011100";
        when "000101111" => n11 <= "0111101011011011";
        when "000110000" => n11 <= "0111101011011010";
        when "000110001" => n11 <= "0111101011011010";
        when "000110010" => n11 <= "0111101011011001";
        when "000110011" => n11 <= "0111100111011000";
        when "000110100" => n11 <= "0111100111010111";
        when "000110101" => n11 <= "0111100111010111";
        when "000110110" => n11 <= "0111100111010110";
        when "000110111" => n11 <= "0111100011010101";
        when "000111000" => n11 <= "0111100011010100";
        when "000111001" => n11 <= "0111100011010100";
        when "000111010" => n11 <= "0111011111010011";
        when "000111011" => n11 <= "0111011111010010";
        when "000111100" => n11 <= "0111011111010001";
        when "000111101" => n11 <= "0111011111010001";
        when "000111110" => n11 <= "0111011011010000";
        when "000111111" => n11 <= "0111011011001111";
        when "001000000" => n11 <= "0111011011001111";
        when "001000001" => n11 <= "0111010111001110";
        when "001000010" => n11 <= "0111010111001101";
        when "001000011" => n11 <= "0111010111001100";
        when "001000100" => n11 <= "0111010111001100";
        when "001000101" => n11 <= "0111010011001011";
        when "001000110" => n11 <= "0111010011001010";
        when "001000111" => n11 <= "0111010011001001";
        when "001001000" => n11 <= "0111001111001001";
        when "001001001" => n11 <= "0111001111001000";
        when "001001010" => n11 <= "0111001111000111";
        when "001001011" => n11 <= "0111001011000111";
        when "001001100" => n11 <= "0111001011000110";
        when "001001101" => n11 <= "0111000111000101";
        when "001001110" => n11 <= "0111000111000101";
        when "001001111" => n11 <= "0111000111000100";
        when "001010000" => n11 <= "0111000011000011";
        when "001010001" => n11 <= "0111000011000010";
        when "001010010" => n11 <= "0111000011000010";
        when "001010011" => n11 <= "0110111111000001";
        when "001010100" => n11 <= "0110111111000000";
        when "001010101" => n11 <= "0110111011000000";
        when "001010110" => n11 <= "0110111010111111";
        when "001010111" => n11 <= "0110111010111110";
        when "001011000" => n11 <= "0110110110111110";
        when "001011001" => n11 <= "0110110110111101";
        when "001011010" => n11 <= "0110110010111100";
        when "001011011" => n11 <= "0110110010111100";
        when "001011100" => n11 <= "0110110010111011";
        when "001011101" => n11 <= "0110101110111010";
        when "001011110" => n11 <= "0110101110111010";
        when "001011111" => n11 <= "0110101010111001";
        when "001100000" => n11 <= "0110101010111000";
        when "001100001" => n11 <= "0110100110111000";
        when "001100010" => n11 <= "0110100110110111";
        when "001100011" => n11 <= "0110100110110110";
        when "001100100" => n11 <= "0110100010110110";
        when "001100101" => n11 <= "0110100010110101";
        when "001100110" => n11 <= "0110011110110101";
        when "001100111" => n11 <= "0110011110110100";
        when "001101000" => n11 <= "0110011010110011";
        when "001101001" => n11 <= "0110011010110011";
        when "001101010" => n11 <= "0110010110110010";
        when "001101011" => n11 <= "0110010110110001";
        when "001101100" => n11 <= "0110010010110001";
        when "001101101" => n11 <= "0110010010110000";
        when "001101110" => n11 <= "0110001110110000";
        when "001101111" => n11 <= "0110001110101111";
        when "001110000" => n11 <= "0110001010101110";
        when "001110001" => n11 <= "0110001010101110";
        when "001110010" => n11 <= "0110000110101101";
        when "001110011" => n11 <= "0110000110101100";
        when "001110100" => n11 <= "0110000010101100";
        when "001110101" => n11 <= "0110000010101011";
        when "001110110" => n11 <= "0101111110101011";
        when "001110111" => n11 <= "0101111110101010";
        when "001111000" => n11 <= "0101111010101010";
        when "001111001" => n11 <= "0101111010101001";
        when "001111010" => n11 <= "0101110110101000";
        when "001111011" => n11 <= "0101110110101000";
        when "001111100" => n11 <= "0101110010100111";
        when "001111101" => n11 <= "0101110010100111";
        when "001111110" => n11 <= "0101101110100110";
        when "001111111" => n11 <= "0101101110100110";
        when "010000000" => n11 <= "0101101010100101";
        when "010000001" => n11 <= "0101100110100100";
        when "010000010" => n11 <= "0101100110100100";
        when "010000011" => n11 <= "0101100010100011";
        when "010000100" => n11 <= "0101100010100011";
        when "010000101" => n11 <= "0101011110100010";
        when "010000110" => n11 <= "0101011110100010";
        when "010000111" => n11 <= "0101011010100001";
        when "010001000" => n11 <= "0101010110100001";
        when "010001001" => n11 <= "0101010110100000";
        when "010001010" => n11 <= "0101010010100000";
        when "010001011" => n11 <= "0101010010011111";
        when "010001100" => n11 <= "0101001110011111";
        when "010001101" => n11 <= "0101001110011110";
        when "010001110" => n11 <= "0101001010011110";
        when "010001111" => n11 <= "0101000110011101";
        when "010010000" => n11 <= "0101000110011101";
        when "010010001" => n11 <= "0101000010011100";
        when "010010010" => n11 <= "0100111110011100";
        when "010010011" => n11 <= "0100111110011011";
        when "010010100" => n11 <= "0100111010011011";
        when "010010101" => n11 <= "0100111010011010";
        when "010010110" => n11 <= "0100110110011010";
        when "010010111" => n11 <= "0100110010011001";
        when "010011000" => n11 <= "0100110010011001";
        when "010011001" => n11 <= "0100101110011000";
        when "010011010" => n11 <= "0100101010011000";
        when "010011011" => n11 <= "0100101010010111";
        when "010011100" => n11 <= "0100100110010111";
        when "010011101" => n11 <= "0100100110010110";
        when "010011110" => n11 <= "0100100010010110";
        when "010011111" => n11 <= "0100011110010110";
        when "010100000" => n11 <= "0100011110010101";
        when "010100001" => n11 <= "0100011010010101";
        when "010100010" => n11 <= "0100010110010100";
        when "010100011" => n11 <= "0100010110010100";
        when "010100100" => n11 <= "0100010010010011";
        when "010100101" => n11 <= "0100001110010011";
        when "010100110" => n11 <= "0100001110010011";
        when "010100111" => n11 <= "0100001010010010";
        when "010101000" => n11 <= "0100000110010010";
        when "010101001" => n11 <= "0100000110010001";
        when "010101010" => n11 <= "0100000010010001";
        when "010101011" => n11 <= "0011111110010001";
        when "010101100" => n11 <= "0011111110010000";
        when "010101101" => n11 <= "0011111010010000";
        when "010101110" => n11 <= "0011110110001111";
        when "010101111" => n11 <= "0011110110001111";
        when "010110000" => n11 <= "0011110010001111";
        when "010110001" => n11 <= "0011101110001110";
        when "010110010" => n11 <= "0011101010001110";
        when "010110011" => n11 <= "0011101010001110";
        when "010110100" => n11 <= "0011100110001101";
        when "010110101" => n11 <= "0011100010001101";
        when "010110110" => n11 <= "0011100010001100";
        when "010110111" => n11 <= "0011011110001100";
        when "010111000" => n11 <= "0011011010001100";
        when "010111001" => n11 <= "0011011010001011";
        when "010111010" => n11 <= "0011010110001011";
        when "010111011" => n11 <= "0011010010001011";
        when "010111100" => n11 <= "0011001110001010";
        when "010111101" => n11 <= "0011001110001010";
        when "010111110" => n11 <= "0011001010001010";
        when "010111111" => n11 <= "0011000110001010";
        when "011000000" => n11 <= "0011000010001001";
        when "011000001" => n11 <= "0011000010001001";
        when "011000010" => n11 <= "0010111110001001";
        when "011000011" => n11 <= "0010111010001000";
        when "011000100" => n11 <= "0010111010001000";
        when "011000101" => n11 <= "0010110110001000";
        when "011000110" => n11 <= "0010110010001000";
        when "011000111" => n11 <= "0010101110000111";
        when "011001000" => n11 <= "0010101110000111";
        when "011001001" => n11 <= "0010101010000111";
        when "011001010" => n11 <= "0010100110000110";
        when "011001011" => n11 <= "0010100010000110";
        when "011001100" => n11 <= "0010100010000110";
        when "011001101" => n11 <= "0010011110000110";
        when "011001110" => n11 <= "0010011010000101";
        when "011001111" => n11 <= "0010010110000101";
        when "011010000" => n11 <= "0010010110000101";
        when "011010001" => n11 <= "0010010010000101";
        when "011010010" => n11 <= "0010001110000101";
        when "011010011" => n11 <= "0010001010000100";
        when "011010100" => n11 <= "0010001010000100";
        when "011010101" => n11 <= "0010000110000100";
        when "011010110" => n11 <= "0010000010000100";
        when "011010111" => n11 <= "0001111110000100";
        when "011011000" => n11 <= "0001111110000011";
        when "011011001" => n11 <= "0001111010000011";
        when "011011010" => n11 <= "0001110110000011";
        when "011011011" => n11 <= "0001110010000011";
        when "011011100" => n11 <= "0001110010000011";
        when "011011101" => n11 <= "0001101110000010";
        when "011011110" => n11 <= "0001101010000010";
        when "011011111" => n11 <= "0001100110000010";
        when "011100000" => n11 <= "0001100010000010";
        when "011100001" => n11 <= "0001100010000010";
        when "011100010" => n11 <= "0001011110000010";
        when "011100011" => n11 <= "0001011010000010";
        when "011100100" => n11 <= "0001010110000001";
        when "011100101" => n11 <= "0001010110000001";
        when "011100110" => n11 <= "0001010010000001";
        when "011100111" => n11 <= "0001001110000001";
        when "011101000" => n11 <= "0001001010000001";
        when "011101001" => n11 <= "0001001010000001";
        when "011101010" => n11 <= "0001000110000001";
        when "011101011" => n11 <= "0001000010000001";
        when "011101100" => n11 <= "0000111110000000";
        when "011101101" => n11 <= "0000111010000000";
        when "011101110" => n11 <= "0000111010000000";
        when "011101111" => n11 <= "0000110110000000";
        when "011110000" => n11 <= "0000110010000000";
        when "011110001" => n11 <= "0000101110000000";
        when "011110010" => n11 <= "0000101010000000";
        when "011110011" => n11 <= "0000101010000000";
        when "011110100" => n11 <= "0000100110000000";
        when "011110101" => n11 <= "0000100010000000";
        when "011110110" => n11 <= "0000011110000000";
        when "011110111" => n11 <= "0000011110000000";
        when "011111000" => n11 <= "0000011010000000";
        when "011111001" => n11 <= "0000010110000000";
        when "011111010" => n11 <= "0000010010000000";
        when "011111011" => n11 <= "0000001110000000";
        when "011111100" => n11 <= "0000001110000000";
        when "011111101" => n11 <= "0000001010000000";
        when "011111110" => n11 <= "0000000110000000";
        when "011111111" => n11 <= "0000000010000000";
        when "100000000" => n11 <= "0000000010000000";
        when "100000001" => n11 <= "1111111110000000";
        when "100000010" => n11 <= "1111111010000000";
        when "100000011" => n11 <= "1111110110000000";
        when "100000100" => n11 <= "1111110010000000";
        when "100000101" => n11 <= "1111110010000000";
        when "100000110" => n11 <= "1111101110000000";
        when "100000111" => n11 <= "1111101010000000";
        when "100001000" => n11 <= "1111100110000000";
        when "100001001" => n11 <= "1111100010000000";
        when "100001010" => n11 <= "1111100010000000";
        when "100001011" => n11 <= "1111011110000000";
        when "100001100" => n11 <= "1111011010000000";
        when "100001101" => n11 <= "1111010110000000";
        when "100001110" => n11 <= "1111010110000000";
        when "100001111" => n11 <= "1111010010000000";
        when "100010000" => n11 <= "1111001110000000";
        when "100010001" => n11 <= "1111001010000000";
        when "100010010" => n11 <= "1111000110000000";
        when "100010011" => n11 <= "1111000110000000";
        when "100010100" => n11 <= "1111000010000000";
        when "100010101" => n11 <= "1110111110000001";
        when "100010110" => n11 <= "1110111010000001";
        when "100010111" => n11 <= "1110110110000001";
        when "100011000" => n11 <= "1110110110000001";
        when "100011001" => n11 <= "1110110010000001";
        when "100011010" => n11 <= "1110101110000001";
        when "100011011" => n11 <= "1110101010000001";
        when "100011100" => n11 <= "1110101010000001";
        when "100011101" => n11 <= "1110100110000010";
        when "100011110" => n11 <= "1110100010000010";
        when "100011111" => n11 <= "1110011110000010";
        when "100100000" => n11 <= "1110011110000010";
        when "100100001" => n11 <= "1110011010000010";
        when "100100010" => n11 <= "1110010110000010";
        when "100100011" => n11 <= "1110010010000010";
        when "100100100" => n11 <= "1110001110000011";
        when "100100101" => n11 <= "1110001110000011";
        when "100100110" => n11 <= "1110001010000011";
        when "100100111" => n11 <= "1110000110000011";
        when "100101000" => n11 <= "1110000010000011";
        when "100101001" => n11 <= "1110000010000100";
        when "100101010" => n11 <= "1101111110000100";
        when "100101011" => n11 <= "1101111010000100";
        when "100101100" => n11 <= "1101110110000100";
        when "100101101" => n11 <= "1101110110000100";
        when "100101110" => n11 <= "1101110010000101";
        when "100101111" => n11 <= "1101101110000101";
        when "100110000" => n11 <= "1101101010000101";
        when "100110001" => n11 <= "1101101010000101";
        when "100110010" => n11 <= "1101100110000101";
        when "100110011" => n11 <= "1101100010000110";
        when "100110100" => n11 <= "1101011110000110";
        when "100110101" => n11 <= "1101011110000110";
        when "100110110" => n11 <= "1101011010000110";
        when "100110111" => n11 <= "1101010110000111";
        when "100111000" => n11 <= "1101010010000111";
        when "100111001" => n11 <= "1101010010000111";
        when "100111010" => n11 <= "1101001110001000";
        when "100111011" => n11 <= "1101001010001000";
        when "100111100" => n11 <= "1101000110001000";
        when "100111101" => n11 <= "1101000110001000";
        when "100111110" => n11 <= "1101000010001001";
        when "100111111" => n11 <= "1100111110001001";
        when "101000000" => n11 <= "1100111110001001";
        when "101000001" => n11 <= "1100111010001010";
        when "101000010" => n11 <= "1100110110001010";
        when "101000011" => n11 <= "1100110010001010";
        when "101000100" => n11 <= "1100110010001010";
        when "101000101" => n11 <= "1100101110001011";
        when "101000110" => n11 <= "1100101010001011";
        when "101000111" => n11 <= "1100100110001011";
        when "101001000" => n11 <= "1100100110001100";
        when "101001001" => n11 <= "1100100010001100";
        when "101001010" => n11 <= "1100011110001100";
        when "101001011" => n11 <= "1100011110001101";
        when "101001100" => n11 <= "1100011010001101";
        when "101001101" => n11 <= "1100010110001110";
        when "101001110" => n11 <= "1100010110001110";
        when "101001111" => n11 <= "1100010010001110";
        when "101010000" => n11 <= "1100001110001111";
        when "101010001" => n11 <= "1100001010001111";
        when "101010010" => n11 <= "1100001010001111";
        when "101010011" => n11 <= "1100000110010000";
        when "101010100" => n11 <= "1100000010010000";
        when "101010101" => n11 <= "1100000010010001";
        when "101010110" => n11 <= "1011111110010001";
        when "101010111" => n11 <= "1011111010010001";
        when "101011000" => n11 <= "1011111010010010";
        when "101011001" => n11 <= "1011110110010010";
        when "101011010" => n11 <= "1011110010010011";
        when "101011011" => n11 <= "1011110010010011";
        when "101011100" => n11 <= "1011101110010011";
        when "101011101" => n11 <= "1011101010010100";
        when "101011110" => n11 <= "1011101010010100";
        when "101011111" => n11 <= "1011100110010101";
        when "101100000" => n11 <= "1011100010010101";
        when "101100001" => n11 <= "1011100010010110";
        when "101100010" => n11 <= "1011011110010110";
        when "101100011" => n11 <= "1011011010010110";
        when "101100100" => n11 <= "1011011010010111";
        when "101100101" => n11 <= "1011010110010111";
        when "101100110" => n11 <= "1011010110011000";
        when "101100111" => n11 <= "1011010010011000";
        when "101101000" => n11 <= "1011001110011001";
        when "101101001" => n11 <= "1011001110011001";
        when "101101010" => n11 <= "1011001010011010";
        when "101101011" => n11 <= "1011000110011010";
        when "101101100" => n11 <= "1011000110011011";
        when "101101101" => n11 <= "1011000010011011";
        when "101101110" => n11 <= "1011000010011100";
        when "101101111" => n11 <= "1010111110011100";
        when "101110000" => n11 <= "1010111010011101";
        when "101110001" => n11 <= "1010111010011101";
        when "101110010" => n11 <= "1010110110011110";
        when "101110011" => n11 <= "1010110010011110";
        when "101110100" => n11 <= "1010110010011111";
        when "101110101" => n11 <= "1010101110011111";
        when "101110110" => n11 <= "1010101110100000";
        when "101110111" => n11 <= "1010101010100000";
        when "101111000" => n11 <= "1010101010100001";
        when "101111001" => n11 <= "1010100110100001";
        when "101111010" => n11 <= "1010100010100010";
        when "101111011" => n11 <= "1010100010100010";
        when "101111100" => n11 <= "1010011110100011";
        when "101111101" => n11 <= "1010011110100011";
        when "101111110" => n11 <= "1010011010100100";
        when "101111111" => n11 <= "1010011010100100";
        when "110000000" => n11 <= "1010010110100101";
        when "110000001" => n11 <= "1010010010100110";
        when "110000010" => n11 <= "1010010010100110";
        when "110000011" => n11 <= "1010001110100111";
        when "110000100" => n11 <= "1010001110100111";
        when "110000101" => n11 <= "1010001010101000";
        when "110000110" => n11 <= "1010001010101000";
        when "110000111" => n11 <= "1010000110101001";
        when "110001000" => n11 <= "1010000110101010";
        when "110001001" => n11 <= "1010000010101010";
        when "110001010" => n11 <= "1010000010101011";
        when "110001011" => n11 <= "1001111110101011";
        when "110001100" => n11 <= "1001111110101100";
        when "110001101" => n11 <= "1001111010101100";
        when "110001110" => n11 <= "1001111010101101";
        when "110001111" => n11 <= "1001110110101110";
        when "110010000" => n11 <= "1001110110101110";
        when "110010001" => n11 <= "1001110010101111";
        when "110010010" => n11 <= "1001110010110000";
        when "110010011" => n11 <= "1001101110110000";
        when "110010100" => n11 <= "1001101110110001";
        when "110010101" => n11 <= "1001101010110001";
        when "110010110" => n11 <= "1001101010110010";
        when "110010111" => n11 <= "1001100110110011";
        when "110011000" => n11 <= "1001100110110011";
        when "110011001" => n11 <= "1001100010110100";
        when "110011010" => n11 <= "1001100010110101";
        when "110011011" => n11 <= "1001011110110101";
        when "110011100" => n11 <= "1001011110110110";
        when "110011101" => n11 <= "1001011010110110";
        when "110011110" => n11 <= "1001011010110111";
        when "110011111" => n11 <= "1001011010111000";
        when "110100000" => n11 <= "1001010110111000";
        when "110100001" => n11 <= "1001010110111001";
        when "110100010" => n11 <= "1001010010111010";
        when "110100011" => n11 <= "1001010010111010";
        when "110100100" => n11 <= "1001001110111011";
        when "110100101" => n11 <= "1001001110111100";
        when "110100110" => n11 <= "1001001110111100";
        when "110100111" => n11 <= "1001001010111101";
        when "110101000" => n11 <= "1001001010111110";
        when "110101001" => n11 <= "1001000110111110";
        when "110101010" => n11 <= "1001000110111111";
        when "110101011" => n11 <= "1001000111000000";
        when "110101100" => n11 <= "1001000011000000";
        when "110101101" => n11 <= "1001000011000001";
        when "110101110" => n11 <= "1000111111000010";
        when "110101111" => n11 <= "1000111111000010";
        when "110110000" => n11 <= "1000111111000011";
        when "110110001" => n11 <= "1000111011000100";
        when "110110010" => n11 <= "1000111011000101";
        when "110110011" => n11 <= "1000111011000101";
        when "110110100" => n11 <= "1000110111000110";
        when "110110101" => n11 <= "1000110111000111";
        when "110110110" => n11 <= "1000110011000111";
        when "110110111" => n11 <= "1000110011001000";
        when "110111000" => n11 <= "1000110011001001";
        when "110111001" => n11 <= "1000101111001001";
        when "110111010" => n11 <= "1000101111001010";
        when "110111011" => n11 <= "1000101111001011";
        when "110111100" => n11 <= "1000101011001100";
        when "110111101" => n11 <= "1000101011001100";
        when "110111110" => n11 <= "1000101011001101";
        when "110111111" => n11 <= "1000101011001110";
        when "111000000" => n11 <= "1000100111001111";
        when "111000001" => n11 <= "1000100111001111";
        when "111000010" => n11 <= "1000100111010000";
        when "111000011" => n11 <= "1000100011010001";
        when "111000100" => n11 <= "1000100011010001";
        when "111000101" => n11 <= "1000100011010010";
        when "111000110" => n11 <= "1000100011010011";
        when "111000111" => n11 <= "1000011111010100";
        when "111001000" => n11 <= "1000011111010100";
        when "111001001" => n11 <= "1000011111010101";
        when "111001010" => n11 <= "1000011011010110";
        when "111001011" => n11 <= "1000011011010111";
        when "111001100" => n11 <= "1000011011010111";
        when "111001101" => n11 <= "1000011011011000";
        when "111001110" => n11 <= "1000010111011001";
        when "111001111" => n11 <= "1000010111011010";
        when "111010000" => n11 <= "1000010111011010";
        when "111010001" => n11 <= "1000010111011011";
        when "111010010" => n11 <= "1000010111011100";
        when "111010011" => n11 <= "1000010011011101";
        when "111010100" => n11 <= "1000010011011101";
        when "111010101" => n11 <= "1000010011011110";
        when "111010110" => n11 <= "1000010011011111";
        when "111010111" => n11 <= "1000010011100000";
        when "111011000" => n11 <= "1000001111100000";
        when "111011001" => n11 <= "1000001111100001";
        when "111011010" => n11 <= "1000001111100010";
        when "111011011" => n11 <= "1000001111100011";
        when "111011100" => n11 <= "1000001111100011";
        when "111011101" => n11 <= "1000001011100100";
        when "111011110" => n11 <= "1000001011100101";
        when "111011111" => n11 <= "1000001011100110";
        when "111100000" => n11 <= "1000001011100111";
        when "111100001" => n11 <= "1000001011100111";
        when "111100010" => n11 <= "1000001011101000";
        when "111100011" => n11 <= "1000001011101001";
        when "111100100" => n11 <= "1000000111101010";
        when "111100101" => n11 <= "1000000111101010";
        when "111100110" => n11 <= "1000000111101011";
        when "111100111" => n11 <= "1000000111101100";
        when "111101000" => n11 <= "1000000111101101";
        when "111101001" => n11 <= "1000000111101101";
        when "111101010" => n11 <= "1000000111101110";
        when "111101011" => n11 <= "1000000111101111";
        when "111101100" => n11 <= "1000000011110000";
        when "111101101" => n11 <= "1000000011110001";
        when "111101110" => n11 <= "1000000011110001";
        when "111101111" => n11 <= "1000000011110010";
        when "111110000" => n11 <= "1000000011110011";
        when "111110001" => n11 <= "1000000011110100";
        when "111110010" => n11 <= "1000000011110101";
        when "111110011" => n11 <= "1000000011110101";
        when "111110100" => n11 <= "1000000011110110";
        when "111110101" => n11 <= "1000000011110111";
        when "111110110" => n11 <= "1000000011111000";
        when "111110111" => n11 <= "1000000011111000";
        when "111111000" => n11 <= "1000000011111001";
        when "111111001" => n11 <= "1000000011111010";
        when "111111010" => n11 <= "1000000011111011";
        when "111111011" => n11 <= "1000000011111100";
        when "111111100" => n11 <= "1000000011111100";
        when "111111101" => n11 <= "1000000011111101";
        when "111111110" => n11 <= "1000000011111110";
        when "111111111" => n11 <= "1000000011111111";
        when others => n11 <= "XXXXXXXXXXXXXXXX";
      end case;
    end if;
  end if;
end process;
n12 <= n11(15 downto 15) &
  n11(14 downto 14) &
  n11(13 downto 13) &
  n11(12 downto 12) &
  n11(11 downto 11) &
  n11(10 downto 10) &
  n11(9 downto 9) &
  n11(8 downto 8);
n13 <= n11(7 downto 7) &
  n11(6 downto 6) &
  n11(5 downto 5) &
  n11(4 downto 4) &
  n11(3 downto 3) &
  n11(2 downto 2) &
  n11(1 downto 1) &
  n11(0 downto 0);
n14 <= unsigned(signed(n5) * signed(n12));
n15 <= n14(14 downto 14) &
  n14(13 downto 13) &
  n14(12 downto 12) &
  n14(11 downto 11) &
  n14(10 downto 10) &
  n14(9 downto 9) &
  n14(8 downto 8) &
  n14(7 downto 7);
process (clock_c) begin
  if rising_edge(clock_c) then
    if i5 = "1" then
      n16 <= "00000000";
    elsif i4 = "1" then
      n16 <= n15;
    end if;
  end if;
end process;
n17 <= unsigned(signed(n6) * signed(n13));
n18 <= n17(14 downto 14) &
  n17(13 downto 13) &
  n17(12 downto 12) &
  n17(11 downto 11) &
  n17(10 downto 10) &
  n17(9 downto 9) &
  n17(8 downto 8) &
  n17(7 downto 7);
process (clock_c) begin
  if rising_edge(clock_c) then
    if i5 = "1" then
      n19 <= "00000000";
    elsif i4 = "1" then
      n19 <= n18;
    end if;
  end if;
end process;
n20 <= n16 - n19;
process (clock_c) begin
  if rising_edge(clock_c) then
    if i5 = "1" then
      n21 <= "00000000";
    elsif i4 = "1" then
      n21 <= n20;
    end if;
  end if;
end process;
n22 <= unsigned(signed(n5) * signed(n13));
n23 <= n22(14 downto 14) &
  n22(13 downto 13) &
  n22(12 downto 12) &
  n22(11 downto 11) &
  n22(10 downto 10) &
  n22(9 downto 9) &
  n22(8 downto 8) &
  n22(7 downto 7);
process (clock_c) begin
  if rising_edge(clock_c) then
    if i5 = "1" then
      n24 <= "00000000";
    elsif i4 = "1" then
      n24 <= n23;
    end if;
  end if;
end process;
n25 <= unsigned(signed(n6) * signed(n12));
n26 <= n25(14 downto 14) &
  n25(13 downto 13) &
  n25(12 downto 12) &
  n25(11 downto 11) &
  n25(10 downto 10) &
  n25(9 downto 9) &
  n25(8 downto 8) &
  n25(7 downto 7);
process (clock_c) begin
  if rising_edge(clock_c) then
    if i5 = "1" then
      n27 <= "00000000";
    elsif i4 = "1" then
      n27 <= n26;
    end if;
  end if;
end process;
n28 <= n24 + n27;
process (clock_c) begin
  if rising_edge(clock_c) then
    if i5 = "1" then
      n29 <= "00000000";
    elsif i4 = "1" then
      n29 <= n28;
    end if;
  end if;
end process;
n30 <= n8 + n21;
n31 <= n10 + n29;
n32 <= n30 & n31;
process (clock_c) begin
  if rising_edge(clock_c) then
    if i5 = "1" then
      n33 <= "0000000000000000";
    elsif i4 = "1" then
      n33 <= n32;
    end if;
  end if;
end process;
n34 <= n8 - n21;
n35 <= n10 - n29;
n36 <= n34 & n35;
process (clock_c) begin
  if rising_edge(clock_c) then
    if i5 = "1" then
      n37 <= "0000000000000000";
    elsif i4 = "1" then
      n37 <= n36;
    end if;
  end if;
end process;
o2 <= n37;
o1 <= n33;
end architecture rtl;

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
entity cf_fft_2048_8_21 is
port (
clock_c : in std_logic;
i1 : in  unsigned(0 downto 0);
i2 : in  unsigned(15 downto 0);
i3 : in  unsigned(15 downto 0);
i4 : in  unsigned(0 downto 0);
i5 : in  unsigned(0 downto 0);
o1 : out unsigned(0 downto 0);
o2 : out unsigned(15 downto 0);
o3 : out unsigned(15 downto 0));
end entity cf_fft_2048_8_21;
architecture rtl of cf_fft_2048_8_21 is
signal n1 : unsigned(8 downto 0);
signal n2 : unsigned(31 downto 0);
signal n3 : unsigned(0 downto 0) := "0";
signal n4 : unsigned(0 downto 0) := "0";
signal n5 : unsigned(0 downto 0) := "0";
signal n6 : unsigned(0 downto 0) := "0";
signal n7 : unsigned(8 downto 0);
signal n8 : unsigned(8 downto 0) := "000000000";
signal n9 : unsigned(8 downto 0) := "000000000";
signal n10 : unsigned(8 downto 0) := "000000000";
signal n11 : unsigned(8 downto 0) := "000000000";
signal n12 : unsigned(0 downto 0);
signal n13 : unsigned(0 downto 0) := "0";
signal n14 : unsigned(0 downto 0) := "0";
signal n15 : unsigned(0 downto 0) := "0";
signal n16 : unsigned(0 downto 0) := "0";
signal n17 : unsigned(0 downto 0);
signal n18 : unsigned(1 downto 0);
signal n19 : unsigned(15 downto 0);
signal n20 : unsigned(15 downto 0);
signal n21 : unsigned(15 downto 0);
signal n22 : unsigned(15 downto 0);
signal n23 : unsigned(15 downto 0);
signal n24 : unsigned(15 downto 0);
signal s25_1 : unsigned(15 downto 0);
signal s25_2 : unsigned(15 downto 0);
signal s26_1 : unsigned(0 downto 0);
signal s27_1 : unsigned(31 downto 0);
signal s28_1 : unsigned(0 downto 0);
signal s28_2 : unsigned(0 downto 0);
signal s28_3 : unsigned(31 downto 0);
signal s29_1 : unsigned(9 downto 0);
signal s29_2 : unsigned(0 downto 0);
component cf_fft_2048_8_22 is
port (
clock_c : in std_logic;
i1 : in  unsigned(15 downto 0);
i2 : in  unsigned(15 downto 0);
i3 : in  unsigned(8 downto 0);
i4 : in  unsigned(0 downto 0);
i5 : in  unsigned(0 downto 0);
o1 : out unsigned(15 downto 0);
o2 : out unsigned(15 downto 0));
end component cf_fft_2048_8_22;
component cf_fft_2048_8_35 is
port (
clock_c : in std_logic;
i1 : in  unsigned(1 downto 0);
i2 : in  unsigned(0 downto 0);
i3 : in  unsigned(0 downto 0);
o1 : out unsigned(0 downto 0));
end component cf_fft_2048_8_35;
component cf_fft_2048_8_31 is
port (
clock_c : in std_logic;
i1 : in  unsigned(31 downto 0);
i2 : in  unsigned(0 downto 0);
i3 : in  unsigned(8 downto 0);
i4 : in  unsigned(0 downto 0);
i5 : in  unsigned(0 downto 0);
i6 : in  unsigned(0 downto 0);
o1 : out unsigned(31 downto 0));
end component cf_fft_2048_8_31;
component cf_fft_2048_8_30 is
port (
clock_c : in std_logic;
i1 : in  unsigned(31 downto 0);
i2 : in  unsigned(0 downto 0);
i3 : in  unsigned(8 downto 0);
i4 : in  unsigned(0 downto 0);
i5 : in  unsigned(0 downto 0);
i6 : in  unsigned(0 downto 0);
o1 : out unsigned(0 downto 0);
o2 : out unsigned(0 downto 0);
o3 : out unsigned(31 downto 0));
end component cf_fft_2048_8_30;
component cf_fft_2048_8_26 is
port (
clock_c : in std_logic;
i1 : in  unsigned(0 downto 0);
i2 : in  unsigned(0 downto 0);
i3 : in  unsigned(0 downto 0);
o1 : out unsigned(9 downto 0);
o2 : out unsigned(0 downto 0));
end component cf_fft_2048_8_26;
begin
n1 <= s29_1(9 downto 9) &
  s29_1(8 downto 8) &
  s29_1(7 downto 7) &
  s29_1(6 downto 6) &
  s29_1(5 downto 5) &
  s29_1(4 downto 4) &
  s29_1(3 downto 3) &
  s29_1(2 downto 2) &
  s29_1(1 downto 1);
n2 <= s25_1 & s25_2;
process (clock_c) begin
  if rising_edge(clock_c) then
    if i5 = "1" then
      n3 <= "0";
    elsif i4 = "1" then
      n3 <= s29_2;
    end if;
  end if;
end process;
process (clock_c) begin
  if rising_edge(clock_c) then
    if i5 = "1" then
      n4 <= "0";
    elsif i4 = "1" then
      n4 <= n3;
    end if;
  end if;
end process;
process (clock_c) begin
  if rising_edge(clock_c) then
    if i5 = "1" then
      n5 <= "0";
    elsif i4 = "1" then
      n5 <= n4;
    end if;
  end if;
end process;
process (clock_c) begin
  if rising_edge(clock_c) then
    if i5 = "1" then
      n6 <= "0";
    elsif i4 = "1" then
      n6 <= n5;
    end if;
  end if;
end process;
n7 <= s29_1(9 downto 9) &
  s29_1(8 downto 8) &
  s29_1(7 downto 7) &
  s29_1(6 downto 6) &
  s29_1(5 downto 5) &
  s29_1(4 downto 4) &
  s29_1(3 downto 3) &
  s29_1(2 downto 2) &
  s29_1(1 downto 1);
process (clock_c) begin
  if rising_edge(clock_c) then
    if i5 = "1" then
      n8 <= "000000000";
    elsif i4 = "1" then
      n8 <= n7;
    end if;
  end if;
end process;
process (clock_c) begin
  if rising_edge(clock_c) then
    if i5 = "1" then
      n9 <= "000000000";
    elsif i4 = "1" then
      n9 <= n8;
    end if;
  end if;
end process;
process (clock_c) begin
  if rising_edge(clock_c) then
    if i5 = "1" then
      n10 <= "000000000";
    elsif i4 = "1" then
      n10 <= n9;
    end if;
  end if;
end process;
process (clock_c) begin
  if rising_edge(clock_c) then
    if i5 = "1" then
      n11 <= "000000000";
    elsif i4 = "1" then
      n11 <= n10;
    end if;
  end if;
end process;
n12 <= s29_1(0 downto 0);
process (clock_c) begin
  if rising_edge(clock_c) then
    if i5 = "1" then
      n13 <= "0";
    elsif i4 = "1" then
      n13 <= n12;
    end if;
  end if;
end process;
process (clock_c) begin
  if rising_edge(clock_c) then
    if i5 = "1" then
      n14 <= "0";
    elsif i4 = "1" then
      n14 <= n13;
    end if;
  end if;
end process;
process (clock_c) begin
  if rising_edge(clock_c) then
    if i5 = "1" then
      n15 <= "0";
    elsif i4 = "1" then
      n15 <= n14;
    end if;
  end if;
end process;
process (clock_c) begin
  if rising_edge(clock_c) then
    if i5 = "1" then
      n16 <= "0";
    elsif i4 = "1" then
      n16 <= n15;
    end if;
  end if;
end process;
n17 <= not n16;
n18 <= s28_2 & s28_1;
n19 <= s28_3(31 downto 31) &
  s28_3(30 downto 30) &
  s28_3(29 downto 29) &
  s28_3(28 downto 28) &
  s28_3(27 downto 27) &
  s28_3(26 downto 26) &
  s28_3(25 downto 25) &
  s28_3(24 downto 24) &
  s28_3(23 downto 23) &
  s28_3(22 downto 22) &
  s28_3(21 downto 21) &
  s28_3(20 downto 20) &
  s28_3(19 downto 19) &
  s28_3(18 downto 18) &
  s28_3(17 downto 17) &
  s28_3(16 downto 16);
n20 <= s28_3(15 downto 15) &
  s28_3(14 downto 14) &
  s28_3(13 downto 13) &
  s28_3(12 downto 12) &
  s28_3(11 downto 11) &
  s28_3(10 downto 10) &
  s28_3(9 downto 9) &
  s28_3(8 downto 8) &
  s28_3(7 downto 7) &
  s28_3(6 downto 6) &
  s28_3(5 downto 5) &
  s28_3(4 downto 4) &
  s28_3(3 downto 3) &
  s28_3(2 downto 2) &
  s28_3(1 downto 1) &
  s28_3(0 downto 0);
n21 <= s27_1(31 downto 31) &
  s27_1(30 downto 30) &
  s27_1(29 downto 29) &
  s27_1(28 downto 28) &
  s27_1(27 downto 27) &
  s27_1(26 downto 26) &
  s27_1(25 downto 25) &
  s27_1(24 downto 24) &
  s27_1(23 downto 23) &
  s27_1(22 downto 22) &
  s27_1(21 downto 21) &
  s27_1(20 downto 20) &
  s27_1(19 downto 19) &
  s27_1(18 downto 18) &
  s27_1(17 downto 17) &
  s27_1(16 downto 16);
n22 <= s27_1(15 downto 15) &
  s27_1(14 downto 14) &
  s27_1(13 downto 13) &
  s27_1(12 downto 12) &
  s27_1(11 downto 11) &
  s27_1(10 downto 10) &
  s27_1(9 downto 9) &
  s27_1(8 downto 8) &
  s27_1(7 downto 7) &
  s27_1(6 downto 6) &
  s27_1(5 downto 5) &
  s27_1(4 downto 4) &
  s27_1(3 downto 3) &
  s27_1(2 downto 2) &
  s27_1(1 downto 1) &
  s27_1(0 downto 0);
n23 <= n20 when s26_1 = "1" else n19;
n24 <= n22 when s26_1 = "1" else n21;
s25 : cf_fft_2048_8_22 port map (clock_c, i2, i3, n1, i4, i5, s25_1, s25_2);
s26 : cf_fft_2048_8_35 port map (clock_c, n18, i4, i5, s26_1);
s27 : cf_fft_2048_8_31 port map (clock_c, n2, n6, n11, n16, i4, i5, s27_1);
s28 : cf_fft_2048_8_30 port map (clock_c, n2, n6, n11, n17, i4, i5, s28_1, s28_2, s28_3);
s29 : cf_fft_2048_8_26 port map (clock_c, i1, i4, i5, s29_1, s29_2);
o3 <= n24;
o2 <= n23;
o1 <= s28_1;
end architecture rtl;

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
entity cf_fft_2048_8_20 is
port (
clock_c : in std_logic;
i1 : in  unsigned(15 downto 0);
i2 : in  unsigned(15 downto 0);
i3 : in  unsigned(7 downto 0);
i4 : in  unsigned(0 downto 0);
i5 : in  unsigned(0 downto 0);
o1 : out unsigned(15 downto 0);
o2 : out unsigned(15 downto 0));
end entity cf_fft_2048_8_20;
architecture rtl of cf_fft_2048_8_20 is
signal n1 : unsigned(15 downto 0) := "0000000000000000";
signal n2 : unsigned(7 downto 0);
signal n3 : unsigned(7 downto 0);
signal n4 : unsigned(15 downto 0) := "0000000000000000";
signal n5 : unsigned(7 downto 0);
signal n6 : unsigned(7 downto 0);
signal n7 : unsigned(7 downto 0) := "00000000";
signal n8 : unsigned(7 downto 0) := "00000000";
signal n9 : unsigned(7 downto 0) := "00000000";
signal n10 : unsigned(7 downto 0) := "00000000";
signal n11 : unsigned(15 downto 0) := "0000000000000000";
signal n12 : unsigned(7 downto 0);
signal n13 : unsigned(7 downto 0);
signal n14 : unsigned(15 downto 0);
signal n15 : unsigned(7 downto 0);
signal n16 : unsigned(7 downto 0) := "00000000";
signal n17 : unsigned(15 downto 0);
signal n18 : unsigned(7 downto 0);
signal n19 : unsigned(7 downto 0) := "00000000";
signal n20 : unsigned(7 downto 0);
signal n21 : unsigned(7 downto 0) := "00000000";
signal n22 : unsigned(15 downto 0);
signal n23 : unsigned(7 downto 0);
signal n24 : unsigned(7 downto 0) := "00000000";
signal n25 : unsigned(15 downto 0);
signal n26 : unsigned(7 downto 0);
signal n27 : unsigned(7 downto 0) := "00000000";
signal n28 : unsigned(7 downto 0);
signal n29 : unsigned(7 downto 0) := "00000000";
signal n30 : unsigned(7 downto 0);
signal n31 : unsigned(7 downto 0);
signal n32 : unsigned(15 downto 0);
signal n33 : unsigned(15 downto 0) := "0000000000000000";
signal n34 : unsigned(7 downto 0);
signal n35 : unsigned(7 downto 0);
signal n36 : unsigned(15 downto 0);
signal n37 : unsigned(15 downto 0) := "0000000000000000";
begin
process (clock_c) begin
  if rising_edge(clock_c) then
    if i5 = "1" then
      n1 <= "0000000000000000";
    elsif i4 = "1" then
      n1 <= i1;
    end if;
  end if;
end process;
n2 <= n1(15 downto 15) &
  n1(14 downto 14) &
  n1(13 downto 13) &
  n1(12 downto 12) &
  n1(11 downto 11) &
  n1(10 downto 10) &
  n1(9 downto 9) &
  n1(8 downto 8);
n3 <= n1(7 downto 7) &
  n1(6 downto 6) &
  n1(5 downto 5) &
  n1(4 downto 4) &
  n1(3 downto 3) &
  n1(2 downto 2) &
  n1(1 downto 1) &
  n1(0 downto 0);
process (clock_c) begin
  if rising_edge(clock_c) then
    if i5 = "1" then
      n4 <= "0000000000000000";
    elsif i4 = "1" then
      n4 <= i2;
    end if;
  end if;
end process;
n5 <= n4(15 downto 15) &
  n4(14 downto 14) &
  n4(13 downto 13) &
  n4(12 downto 12) &
  n4(11 downto 11) &
  n4(10 downto 10) &
  n4(9 downto 9) &
  n4(8 downto 8);
n6 <= n4(7 downto 7) &
  n4(6 downto 6) &
  n4(5 downto 5) &
  n4(4 downto 4) &
  n4(3 downto 3) &
  n4(2 downto 2) &
  n4(1 downto 1) &
  n4(0 downto 0);
process (clock_c) begin
  if rising_edge(clock_c) then
    if i5 = "1" then
      n7 <= "00000000";
    elsif i4 = "1" then
      n7 <= n2;
    end if;
  end if;
end process;
process (clock_c) begin
  if rising_edge(clock_c) then
    if i5 = "1" then
      n8 <= "00000000";
    elsif i4 = "1" then
      n8 <= n7;
    end if;
  end if;
end process;
process (clock_c) begin
  if rising_edge(clock_c) then
    if i5 = "1" then
      n9 <= "00000000";
    elsif i4 = "1" then
      n9 <= n3;
    end if;
  end if;
end process;
process (clock_c) begin
  if rising_edge(clock_c) then
    if i5 = "1" then
      n10 <= "00000000";
    elsif i4 = "1" then
      n10 <= n9;
    end if;
  end if;
end process;
process (clock_c) begin
  if rising_edge(clock_c) then 
    if i4 = "1" then
      case i3 is
        when "00000000" => n11 <= "0111111100000000";
        when "00000001" => n11 <= "0111111111111110";
        when "00000010" => n11 <= "0111111111111100";
        when "00000011" => n11 <= "0111111111111011";
        when "00000100" => n11 <= "0111111111111001";
        when "00000101" => n11 <= "0111111111111000";
        when "00000110" => n11 <= "0111111111110110";
        when "00000111" => n11 <= "0111111111110101";
        when "00001000" => n11 <= "0111111111110011";
        when "00001001" => n11 <= "0111111111110001";
        when "00001010" => n11 <= "0111111111110000";
        when "00001011" => n11 <= "0111111011101110";
        when "00001100" => n11 <= "0111111011101101";
        when "00001101" => n11 <= "0111111011101011";
        when "00001110" => n11 <= "0111111011101010";
        when "00001111" => n11 <= "0111110111101000";
        when "00010000" => n11 <= "0111110111100111";
        when "00010001" => n11 <= "0111110111100101";
        when "00010010" => n11 <= "0111110011100011";
        when "00010011" => n11 <= "0111110011100010";
        when "00010100" => n11 <= "0111110011100000";
        when "00010101" => n11 <= "0111101111011111";
        when "00010110" => n11 <= "0111101111011101";
        when "00010111" => n11 <= "0111101011011100";
        when "00011000" => n11 <= "0111101011011010";
        when "00011001" => n11 <= "0111101011011001";
        when "00011010" => n11 <= "0111100111010111";
        when "00011011" => n11 <= "0111100111010110";
        when "00011100" => n11 <= "0111100011010100";
        when "00011101" => n11 <= "0111011111010011";
        when "00011110" => n11 <= "0111011111010001";
        when "00011111" => n11 <= "0111011011010000";
        when "00100000" => n11 <= "0111011011001111";
        when "00100001" => n11 <= "0111010111001101";
        when "00100010" => n11 <= "0111010111001100";
        when "00100011" => n11 <= "0111010011001010";
        when "00100100" => n11 <= "0111001111001001";
        when "00100101" => n11 <= "0111001111000111";
        when "00100110" => n11 <= "0111001011000110";
        when "00100111" => n11 <= "0111000111000101";
        when "00101000" => n11 <= "0111000011000011";
        when "00101001" => n11 <= "0111000011000010";
        when "00101010" => n11 <= "0110111111000000";
        when "00101011" => n11 <= "0110111010111111";
        when "00101100" => n11 <= "0110110110111110";
        when "00101101" => n11 <= "0110110010111100";
        when "00101110" => n11 <= "0110110010111011";
        when "00101111" => n11 <= "0110101110111010";
        when "00110000" => n11 <= "0110101010111000";
        when "00110001" => n11 <= "0110100110110111";
        when "00110010" => n11 <= "0110100010110110";
        when "00110011" => n11 <= "0110011110110101";
        when "00110100" => n11 <= "0110011010110011";
        when "00110101" => n11 <= "0110010110110010";
        when "00110110" => n11 <= "0110010010110001";
        when "00110111" => n11 <= "0110001110110000";
        when "00111000" => n11 <= "0110001010101110";
        when "00111001" => n11 <= "0110000110101101";
        when "00111010" => n11 <= "0110000010101100";
        when "00111011" => n11 <= "0101111110101011";
        when "00111100" => n11 <= "0101111010101010";
        when "00111101" => n11 <= "0101110110101000";
        when "00111110" => n11 <= "0101110010100111";
        when "00111111" => n11 <= "0101101110100110";
        when "01000000" => n11 <= "0101101010100101";
        when "01000001" => n11 <= "0101100110100100";
        when "01000010" => n11 <= "0101100010100011";
        when "01000011" => n11 <= "0101011110100010";
        when "01000100" => n11 <= "0101010110100001";
        when "01000101" => n11 <= "0101010010100000";
        when "01000110" => n11 <= "0101001110011111";
        when "01000111" => n11 <= "0101001010011110";
        when "01001000" => n11 <= "0101000110011101";
        when "01001001" => n11 <= "0100111110011100";
        when "01001010" => n11 <= "0100111010011011";
        when "01001011" => n11 <= "0100110110011010";
        when "01001100" => n11 <= "0100110010011001";
        when "01001101" => n11 <= "0100101010011000";
        when "01001110" => n11 <= "0100100110010111";
        when "01001111" => n11 <= "0100100010010110";
        when "01010000" => n11 <= "0100011110010101";
        when "01010001" => n11 <= "0100010110010100";
        when "01010010" => n11 <= "0100010010010011";
        when "01010011" => n11 <= "0100001110010011";
        when "01010100" => n11 <= "0100000110010010";
        when "01010101" => n11 <= "0100000010010001";
        when "01010110" => n11 <= "0011111110010000";
        when "01010111" => n11 <= "0011110110001111";
        when "01011000" => n11 <= "0011110010001111";
        when "01011001" => n11 <= "0011101010001110";
        when "01011010" => n11 <= "0011100110001101";
        when "01011011" => n11 <= "0011100010001100";
        when "01011100" => n11 <= "0011011010001100";
        when "01011101" => n11 <= "0011010110001011";
        when "01011110" => n11 <= "0011001110001010";
        when "01011111" => n11 <= "0011001010001010";
        when "01100000" => n11 <= "0011000010001001";
        when "01100001" => n11 <= "0010111110001001";
        when "01100010" => n11 <= "0010111010001000";
        when "01100011" => n11 <= "0010110010001000";
        when "01100100" => n11 <= "0010101110000111";
        when "01100101" => n11 <= "0010100110000110";
        when "01100110" => n11 <= "0010100010000110";
        when "01100111" => n11 <= "0010011010000101";
        when "01101000" => n11 <= "0010010110000101";
        when "01101001" => n11 <= "0010001110000101";
        when "01101010" => n11 <= "0010001010000100";
        when "01101011" => n11 <= "0010000010000100";
        when "01101100" => n11 <= "0001111110000011";
        when "01101101" => n11 <= "0001110110000011";
        when "01101110" => n11 <= "0001110010000011";
        when "01101111" => n11 <= "0001101010000010";
        when "01110000" => n11 <= "0001100010000010";
        when "01110001" => n11 <= "0001011110000010";
        when "01110010" => n11 <= "0001010110000001";
        when "01110011" => n11 <= "0001010010000001";
        when "01110100" => n11 <= "0001001010000001";
        when "01110101" => n11 <= "0001000110000001";
        when "01110110" => n11 <= "0000111110000000";
        when "01110111" => n11 <= "0000111010000000";
        when "01111000" => n11 <= "0000110010000000";
        when "01111001" => n11 <= "0000101010000000";
        when "01111010" => n11 <= "0000100110000000";
        when "01111011" => n11 <= "0000011110000000";
        when "01111100" => n11 <= "0000011010000000";
        when "01111101" => n11 <= "0000010010000000";
        when "01111110" => n11 <= "0000001110000000";
        when "01111111" => n11 <= "0000000110000000";
        when "10000000" => n11 <= "0000000010000000";
        when "10000001" => n11 <= "1111111010000000";
        when "10000010" => n11 <= "1111110010000000";
        when "10000011" => n11 <= "1111101110000000";
        when "10000100" => n11 <= "1111100110000000";
        when "10000101" => n11 <= "1111100010000000";
        when "10000110" => n11 <= "1111011010000000";
        when "10000111" => n11 <= "1111010110000000";
        when "10001000" => n11 <= "1111001110000000";
        when "10001001" => n11 <= "1111000110000000";
        when "10001010" => n11 <= "1111000010000000";
        when "10001011" => n11 <= "1110111010000001";
        when "10001100" => n11 <= "1110110110000001";
        when "10001101" => n11 <= "1110101110000001";
        when "10001110" => n11 <= "1110101010000001";
        when "10001111" => n11 <= "1110100010000010";
        when "10010000" => n11 <= "1110011110000010";
        when "10010001" => n11 <= "1110010110000010";
        when "10010010" => n11 <= "1110001110000011";
        when "10010011" => n11 <= "1110001010000011";
        when "10010100" => n11 <= "1110000010000011";
        when "10010101" => n11 <= "1101111110000100";
        when "10010110" => n11 <= "1101110110000100";
        when "10010111" => n11 <= "1101110010000101";
        when "10011000" => n11 <= "1101101010000101";
        when "10011001" => n11 <= "1101100110000101";
        when "10011010" => n11 <= "1101011110000110";
        when "10011011" => n11 <= "1101011010000110";
        when "10011100" => n11 <= "1101010010000111";
        when "10011101" => n11 <= "1101001110001000";
        when "10011110" => n11 <= "1101000110001000";
        when "10011111" => n11 <= "1101000010001001";
        when "10100000" => n11 <= "1100111110001001";
        when "10100001" => n11 <= "1100110110001010";
        when "10100010" => n11 <= "1100110010001010";
        when "10100011" => n11 <= "1100101010001011";
        when "10100100" => n11 <= "1100100110001100";
        when "10100101" => n11 <= "1100011110001100";
        when "10100110" => n11 <= "1100011010001101";
        when "10100111" => n11 <= "1100010110001110";
        when "10101000" => n11 <= "1100001110001111";
        when "10101001" => n11 <= "1100001010001111";
        when "10101010" => n11 <= "1100000010010000";
        when "10101011" => n11 <= "1011111110010001";
        when "10101100" => n11 <= "1011111010010010";
        when "10101101" => n11 <= "1011110010010011";
        when "10101110" => n11 <= "1011101110010011";
        when "10101111" => n11 <= "1011101010010100";
        when "10110000" => n11 <= "1011100010010101";
        when "10110001" => n11 <= "1011011110010110";
        when "10110010" => n11 <= "1011011010010111";
        when "10110011" => n11 <= "1011010110011000";
        when "10110100" => n11 <= "1011001110011001";
        when "10110101" => n11 <= "1011001010011010";
        when "10110110" => n11 <= "1011000110011011";
        when "10110111" => n11 <= "1011000010011100";
        when "10111000" => n11 <= "1010111010011101";
        when "10111001" => n11 <= "1010110110011110";
        when "10111010" => n11 <= "1010110010011111";
        when "10111011" => n11 <= "1010101110100000";
        when "10111100" => n11 <= "1010101010100001";
        when "10111101" => n11 <= "1010100010100010";
        when "10111110" => n11 <= "1010011110100011";
        when "10111111" => n11 <= "1010011010100100";
        when "11000000" => n11 <= "1010010110100101";
        when "11000001" => n11 <= "1010010010100110";
        when "11000010" => n11 <= "1010001110100111";
        when "11000011" => n11 <= "1010001010101000";
        when "11000100" => n11 <= "1010000110101010";
        when "11000101" => n11 <= "1010000010101011";
        when "11000110" => n11 <= "1001111110101100";
        when "11000111" => n11 <= "1001111010101101";
        when "11001000" => n11 <= "1001110110101110";
        when "11001001" => n11 <= "1001110010110000";
        when "11001010" => n11 <= "1001101110110001";
        when "11001011" => n11 <= "1001101010110010";
        when "11001100" => n11 <= "1001100110110011";
        when "11001101" => n11 <= "1001100010110101";
        when "11001110" => n11 <= "1001011110110110";
        when "11001111" => n11 <= "1001011010110111";
        when "11010000" => n11 <= "1001010110111000";
        when "11010001" => n11 <= "1001010010111010";
        when "11010010" => n11 <= "1001001110111011";
        when "11010011" => n11 <= "1001001110111100";
        when "11010100" => n11 <= "1001001010111110";
        when "11010101" => n11 <= "1001000110111111";
        when "11010110" => n11 <= "1001000011000000";
        when "11010111" => n11 <= "1000111111000010";
        when "11011000" => n11 <= "1000111111000011";
        when "11011001" => n11 <= "1000111011000101";
        when "11011010" => n11 <= "1000110111000110";
        when "11011011" => n11 <= "1000110011000111";
        when "11011100" => n11 <= "1000110011001001";
        when "11011101" => n11 <= "1000101111001010";
        when "11011110" => n11 <= "1000101011001100";
        when "11011111" => n11 <= "1000101011001101";
        when "11100000" => n11 <= "1000100111001111";
        when "11100001" => n11 <= "1000100111010000";
        when "11100010" => n11 <= "1000100011010001";
        when "11100011" => n11 <= "1000100011010011";
        when "11100100" => n11 <= "1000011111010100";
        when "11100101" => n11 <= "1000011011010110";
        when "11100110" => n11 <= "1000011011010111";
        when "11100111" => n11 <= "1000010111011001";
        when "11101000" => n11 <= "1000010111011010";
        when "11101001" => n11 <= "1000010111011100";
        when "11101010" => n11 <= "1000010011011101";
        when "11101011" => n11 <= "1000010011011111";
        when "11101100" => n11 <= "1000001111100000";
        when "11101101" => n11 <= "1000001111100010";
        when "11101110" => n11 <= "1000001111100011";
        when "11101111" => n11 <= "1000001011100101";
        when "11110000" => n11 <= "1000001011100111";
        when "11110001" => n11 <= "1000001011101000";
        when "11110010" => n11 <= "1000000111101010";
        when "11110011" => n11 <= "1000000111101011";
        when "11110100" => n11 <= "1000000111101101";
        when "11110101" => n11 <= "1000000111101110";
        when "11110110" => n11 <= "1000000011110000";
        when "11110111" => n11 <= "1000000011110001";
        when "11111000" => n11 <= "1000000011110011";
        when "11111001" => n11 <= "1000000011110101";
        when "11111010" => n11 <= "1000000011110110";
        when "11111011" => n11 <= "1000000011111000";
        when "11111100" => n11 <= "1000000011111001";
        when "11111101" => n11 <= "1000000011111011";
        when "11111110" => n11 <= "1000000011111100";
        when "11111111" => n11 <= "1000000011111110";
        when others => n11 <= "XXXXXXXXXXXXXXXX";
      end case;
    end if;
  end if;
end process;
n12 <= n11(15 downto 15) &
  n11(14 downto 14) &
  n11(13 downto 13) &
  n11(12 downto 12) &
  n11(11 downto 11) &
  n11(10 downto 10) &
  n11(9 downto 9) &
  n11(8 downto 8);
n13 <= n11(7 downto 7) &
  n11(6 downto 6) &
  n11(5 downto 5) &
  n11(4 downto 4) &
  n11(3 downto 3) &
  n11(2 downto 2) &
  n11(1 downto 1) &
  n11(0 downto 0);
n14 <= unsigned(signed(n5) * signed(n12));
n15 <= n14(14 downto 14) &
  n14(13 downto 13) &
  n14(12 downto 12) &
  n14(11 downto 11) &
  n14(10 downto 10) &
  n14(9 downto 9) &
  n14(8 downto 8) &
  n14(7 downto 7);
process (clock_c) begin
  if rising_edge(clock_c) then
    if i5 = "1" then
      n16 <= "00000000";
    elsif i4 = "1" then
      n16 <= n15;
    end if;
  end if;
end process;
n17 <= unsigned(signed(n6) * signed(n13));
n18 <= n17(14 downto 14) &
  n17(13 downto 13) &
  n17(12 downto 12) &
  n17(11 downto 11) &
  n17(10 downto 10) &
  n17(9 downto 9) &
  n17(8 downto 8) &
  n17(7 downto 7);
process (clock_c) begin
  if rising_edge(clock_c) then
    if i5 = "1" then
      n19 <= "00000000";
    elsif i4 = "1" then
      n19 <= n18;
    end if;
  end if;
end process;
n20 <= n16 - n19;
process (clock_c) begin
  if rising_edge(clock_c) then
    if i5 = "1" then
      n21 <= "00000000";
    elsif i4 = "1" then
      n21 <= n20;
    end if;
  end if;
end process;
n22 <= unsigned(signed(n5) * signed(n13));
n23 <= n22(14 downto 14) &
  n22(13 downto 13) &
  n22(12 downto 12) &
  n22(11 downto 11) &
  n22(10 downto 10) &
  n22(9 downto 9) &
  n22(8 downto 8) &
  n22(7 downto 7);
process (clock_c) begin
  if rising_edge(clock_c) then
    if i5 = "1" then
      n24 <= "00000000";
    elsif i4 = "1" then
      n24 <= n23;
    end if;
  end if;
end process;
n25 <= unsigned(signed(n6) * signed(n12));
n26 <= n25(14 downto 14) &
  n25(13 downto 13) &
  n25(12 downto 12) &
  n25(11 downto 11) &
  n25(10 downto 10) &
  n25(9 downto 9) &
  n25(8 downto 8) &
  n25(7 downto 7);
process (clock_c) begin
  if rising_edge(clock_c) then
    if i5 = "1" then
      n27 <= "00000000";
    elsif i4 = "1" then
      n27 <= n26;
    end if;
  end if;
end process;
n28 <= n24 + n27;
process (clock_c) begin
  if rising_edge(clock_c) then
    if i5 = "1" then
      n29 <= "00000000";
    elsif i4 = "1" then
      n29 <= n28;
    end if;
  end if;
end process;
n30 <= n8 + n21;
n31 <= n10 + n29;
n32 <= n30 & n31;
process (clock_c) begin
  if rising_edge(clock_c) then
    if i5 = "1" then
      n33 <= "0000000000000000";
    elsif i4 = "1" then
      n33 <= n32;
    end if;
  end if;
end process;
n34 <= n8 - n21;
n35 <= n10 - n29;
n36 <= n34 & n35;
process (clock_c) begin
  if rising_edge(clock_c) then
    if i5 = "1" then
      n37 <= "0000000000000000";
    elsif i4 = "1" then
      n37 <= n36;
    end if;
  end if;
end process;
o2 <= n37;
o1 <= n33;
end architecture rtl;

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
entity cf_fft_2048_8_19 is
port (
clock_c : in std_logic;
i1 : in  unsigned(0 downto 0);
i2 : in  unsigned(15 downto 0);
i3 : in  unsigned(15 downto 0);
i4 : in  unsigned(0 downto 0);
i5 : in  unsigned(0 downto 0);
o1 : out unsigned(0 downto 0);
o2 : out unsigned(15 downto 0);
o3 : out unsigned(15 downto 0));
end entity cf_fft_2048_8_19;
architecture rtl of cf_fft_2048_8_19 is
signal n1 : unsigned(7 downto 0);
signal n2 : unsigned(31 downto 0);
signal n3 : unsigned(0 downto 0) := "0";
signal n4 : unsigned(0 downto 0) := "0";
signal n5 : unsigned(0 downto 0) := "0";
signal n6 : unsigned(0 downto 0) := "0";
signal n7 : unsigned(8 downto 0);
signal n8 : unsigned(8 downto 0) := "000000000";
signal n9 : unsigned(8 downto 0) := "000000000";
signal n10 : unsigned(8 downto 0) := "000000000";
signal n11 : unsigned(8 downto 0) := "000000000";
signal n12 : unsigned(0 downto 0);
signal n13 : unsigned(0 downto 0) := "0";
signal n14 : unsigned(0 downto 0) := "0";
signal n15 : unsigned(0 downto 0) := "0";
signal n16 : unsigned(0 downto 0) := "0";
signal n17 : unsigned(0 downto 0);
signal n18 : unsigned(1 downto 0);
signal n19 : unsigned(15 downto 0);
signal n20 : unsigned(15 downto 0);
signal n21 : unsigned(15 downto 0);
signal n22 : unsigned(15 downto 0);
signal n23 : unsigned(15 downto 0);
signal n24 : unsigned(15 downto 0);
signal s25_1 : unsigned(15 downto 0);
signal s25_2 : unsigned(15 downto 0);
signal s26_1 : unsigned(0 downto 0);
signal s27_1 : unsigned(31 downto 0);
signal s28_1 : unsigned(0 downto 0);
signal s28_2 : unsigned(0 downto 0);
signal s28_3 : unsigned(31 downto 0);
signal s29_1 : unsigned(9 downto 0);
signal s29_2 : unsigned(0 downto 0);
component cf_fft_2048_8_20 is
port (
clock_c : in std_logic;
i1 : in  unsigned(15 downto 0);
i2 : in  unsigned(15 downto 0);
i3 : in  unsigned(7 downto 0);
i4 : in  unsigned(0 downto 0);
i5 : in  unsigned(0 downto 0);
o1 : out unsigned(15 downto 0);
o2 : out unsigned(15 downto 0));
end component cf_fft_2048_8_20;
component cf_fft_2048_8_35 is
port (
clock_c : in std_logic;
i1 : in  unsigned(1 downto 0);
i2 : in  unsigned(0 downto 0);
i3 : in  unsigned(0 downto 0);
o1 : out unsigned(0 downto 0));
end component cf_fft_2048_8_35;
component cf_fft_2048_8_31 is
port (
clock_c : in std_logic;
i1 : in  unsigned(31 downto 0);
i2 : in  unsigned(0 downto 0);
i3 : in  unsigned(8 downto 0);
i4 : in  unsigned(0 downto 0);
i5 : in  unsigned(0 downto 0);
i6 : in  unsigned(0 downto 0);
o1 : out unsigned(31 downto 0));
end component cf_fft_2048_8_31;
component cf_fft_2048_8_30 is
port (
clock_c : in std_logic;
i1 : in  unsigned(31 downto 0);
i2 : in  unsigned(0 downto 0);
i3 : in  unsigned(8 downto 0);
i4 : in  unsigned(0 downto 0);
i5 : in  unsigned(0 downto 0);
i6 : in  unsigned(0 downto 0);
o1 : out unsigned(0 downto 0);
o2 : out unsigned(0 downto 0);
o3 : out unsigned(31 downto 0));
end component cf_fft_2048_8_30;
component cf_fft_2048_8_26 is
port (
clock_c : in std_logic;
i1 : in  unsigned(0 downto 0);
i2 : in  unsigned(0 downto 0);
i3 : in  unsigned(0 downto 0);
o1 : out unsigned(9 downto 0);
o2 : out unsigned(0 downto 0));
end component cf_fft_2048_8_26;
begin
n1 <= s29_1(9 downto 9) &
  s29_1(8 downto 8) &
  s29_1(7 downto 7) &
  s29_1(6 downto 6) &
  s29_1(5 downto 5) &
  s29_1(4 downto 4) &
  s29_1(3 downto 3) &
  s29_1(2 downto 2);
n2 <= s25_1 & s25_2;
process (clock_c) begin
  if rising_edge(clock_c) then
    if i5 = "1" then
      n3 <= "0";
    elsif i4 = "1" then
      n3 <= s29_2;
    end if;
  end if;
end process;
process (clock_c) begin
  if rising_edge(clock_c) then
    if i5 = "1" then
      n4 <= "0";
    elsif i4 = "1" then
      n4 <= n3;
    end if;
  end if;
end process;
process (clock_c) begin
  if rising_edge(clock_c) then
    if i5 = "1" then
      n5 <= "0";
    elsif i4 = "1" then
      n5 <= n4;
    end if;
  end if;
end process;
process (clock_c) begin
  if rising_edge(clock_c) then
    if i5 = "1" then
      n6 <= "0";
    elsif i4 = "1" then
      n6 <= n5;
    end if;
  end if;
end process;
n7 <= s29_1(9 downto 9) &
  s29_1(8 downto 8) &
  s29_1(7 downto 7) &
  s29_1(6 downto 6) &
  s29_1(5 downto 5) &
  s29_1(4 downto 4) &
  s29_1(3 downto 3) &
  s29_1(2 downto 2) &
  s29_1(1 downto 1);
process (clock_c) begin
  if rising_edge(clock_c) then
    if i5 = "1" then
      n8 <= "000000000";
    elsif i4 = "1" then
      n8 <= n7;
    end if;
  end if;
end process;
process (clock_c) begin
  if rising_edge(clock_c) then
    if i5 = "1" then
      n9 <= "000000000";
    elsif i4 = "1" then
      n9 <= n8;
    end if;
  end if;
end process;
process (clock_c) begin
  if rising_edge(clock_c) then
    if i5 = "1" then
      n10 <= "000000000";
    elsif i4 = "1" then
      n10 <= n9;
    end if;
  end if;
end process;
process (clock_c) begin
  if rising_edge(clock_c) then
    if i5 = "1" then
      n11 <= "000000000";
    elsif i4 = "1" then
      n11 <= n10;
    end if;
  end if;
end process;
n12 <= s29_1(0 downto 0);
process (clock_c) begin
  if rising_edge(clock_c) then
    if i5 = "1" then
      n13 <= "0";
    elsif i4 = "1" then
      n13 <= n12;
    end if;
  end if;
end process;
process (clock_c) begin
  if rising_edge(clock_c) then
    if i5 = "1" then
      n14 <= "0";
    elsif i4 = "1" then
      n14 <= n13;
    end if;
  end if;
end process;
process (clock_c) begin
  if rising_edge(clock_c) then
    if i5 = "1" then
      n15 <= "0";
    elsif i4 = "1" then
      n15 <= n14;
    end if;
  end if;
end process;
process (clock_c) begin
  if rising_edge(clock_c) then
    if i5 = "1" then
      n16 <= "0";
    elsif i4 = "1" then
      n16 <= n15;
    end if;
  end if;
end process;
n17 <= not n16;
n18 <= s28_2 & s28_1;
n19 <= s28_3(31 downto 31) &
  s28_3(30 downto 30) &
  s28_3(29 downto 29) &
  s28_3(28 downto 28) &
  s28_3(27 downto 27) &
  s28_3(26 downto 26) &
  s28_3(25 downto 25) &
  s28_3(24 downto 24) &
  s28_3(23 downto 23) &
  s28_3(22 downto 22) &
  s28_3(21 downto 21) &
  s28_3(20 downto 20) &
  s28_3(19 downto 19) &
  s28_3(18 downto 18) &
  s28_3(17 downto 17) &
  s28_3(16 downto 16);
n20 <= s28_3(15 downto 15) &
  s28_3(14 downto 14) &
  s28_3(13 downto 13) &
  s28_3(12 downto 12) &
  s28_3(11 downto 11) &
  s28_3(10 downto 10) &
  s28_3(9 downto 9) &
  s28_3(8 downto 8) &
  s28_3(7 downto 7) &
  s28_3(6 downto 6) &
  s28_3(5 downto 5) &
  s28_3(4 downto 4) &
  s28_3(3 downto 3) &
  s28_3(2 downto 2) &
  s28_3(1 downto 1) &
  s28_3(0 downto 0);
n21 <= s27_1(31 downto 31) &
  s27_1(30 downto 30) &
  s27_1(29 downto 29) &
  s27_1(28 downto 28) &
  s27_1(27 downto 27) &
  s27_1(26 downto 26) &
  s27_1(25 downto 25) &
  s27_1(24 downto 24) &
  s27_1(23 downto 23) &
  s27_1(22 downto 22) &
  s27_1(21 downto 21) &
  s27_1(20 downto 20) &
  s27_1(19 downto 19) &
  s27_1(18 downto 18) &
  s27_1(17 downto 17) &
  s27_1(16 downto 16);
n22 <= s27_1(15 downto 15) &
  s27_1(14 downto 14) &
  s27_1(13 downto 13) &
  s27_1(12 downto 12) &
  s27_1(11 downto 11) &
  s27_1(10 downto 10) &
  s27_1(9 downto 9) &
  s27_1(8 downto 8) &
  s27_1(7 downto 7) &
  s27_1(6 downto 6) &
  s27_1(5 downto 5) &
  s27_1(4 downto 4) &
  s27_1(3 downto 3) &
  s27_1(2 downto 2) &
  s27_1(1 downto 1) &
  s27_1(0 downto 0);
n23 <= n20 when s26_1 = "1" else n19;
n24 <= n22 when s26_1 = "1" else n21;
s25 : cf_fft_2048_8_20 port map (clock_c, i2, i3, n1, i4, i5, s25_1, s25_2);
s26 : cf_fft_2048_8_35 port map (clock_c, n18, i4, i5, s26_1);
s27 : cf_fft_2048_8_31 port map (clock_c, n2, n6, n11, n16, i4, i5, s27_1);
s28 : cf_fft_2048_8_30 port map (clock_c, n2, n6, n11, n17, i4, i5, s28_1, s28_2, s28_3);
s29 : cf_fft_2048_8_26 port map (clock_c, i1, i4, i5, s29_1, s29_2);
o3 <= n24;
o2 <= n23;
o1 <= s28_1;
end architecture rtl;

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
entity cf_fft_2048_8_18 is
port (
clock_c : in std_logic;
i1 : in  unsigned(15 downto 0);
i2 : in  unsigned(15 downto 0);
i3 : in  unsigned(6 downto 0);
i4 : in  unsigned(0 downto 0);
i5 : in  unsigned(0 downto 0);
o1 : out unsigned(15 downto 0);
o2 : out unsigned(15 downto 0));
end entity cf_fft_2048_8_18;
architecture rtl of cf_fft_2048_8_18 is
signal n1 : unsigned(15 downto 0) := "0000000000000000";
signal n2 : unsigned(7 downto 0);
signal n3 : unsigned(7 downto 0);
signal n4 : unsigned(15 downto 0) := "0000000000000000";
signal n5 : unsigned(7 downto 0);
signal n6 : unsigned(7 downto 0);
signal n7 : unsigned(7 downto 0) := "00000000";
signal n8 : unsigned(7 downto 0) := "00000000";
signal n9 : unsigned(7 downto 0) := "00000000";
signal n10 : unsigned(7 downto 0) := "00000000";
signal n11 : unsigned(15 downto 0) := "0000000000000000";
signal n12 : unsigned(7 downto 0);
signal n13 : unsigned(7 downto 0);
signal n14 : unsigned(15 downto 0);
signal n15 : unsigned(7 downto 0);
signal n16 : unsigned(7 downto 0) := "00000000";
signal n17 : unsigned(15 downto 0);
signal n18 : unsigned(7 downto 0);
signal n19 : unsigned(7 downto 0) := "00000000";
signal n20 : unsigned(7 downto 0);
signal n21 : unsigned(7 downto 0) := "00000000";
signal n22 : unsigned(15 downto 0);
signal n23 : unsigned(7 downto 0);
signal n24 : unsigned(7 downto 0) := "00000000";
signal n25 : unsigned(15 downto 0);
signal n26 : unsigned(7 downto 0);
signal n27 : unsigned(7 downto 0) := "00000000";
signal n28 : unsigned(7 downto 0);
signal n29 : unsigned(7 downto 0) := "00000000";
signal n30 : unsigned(7 downto 0);
signal n31 : unsigned(7 downto 0);
signal n32 : unsigned(15 downto 0);
signal n33 : unsigned(15 downto 0) := "0000000000000000";
signal n34 : unsigned(7 downto 0);
signal n35 : unsigned(7 downto 0);
signal n36 : unsigned(15 downto 0);
signal n37 : unsigned(15 downto 0) := "0000000000000000";
begin
process (clock_c) begin
  if rising_edge(clock_c) then
    if i5 = "1" then
      n1 <= "0000000000000000";
    elsif i4 = "1" then
      n1 <= i1;
    end if;
  end if;
end process;
n2 <= n1(15 downto 15) &
  n1(14 downto 14) &
  n1(13 downto 13) &
  n1(12 downto 12) &
  n1(11 downto 11) &
  n1(10 downto 10) &
  n1(9 downto 9) &
  n1(8 downto 8);
n3 <= n1(7 downto 7) &
  n1(6 downto 6) &
  n1(5 downto 5) &
  n1(4 downto 4) &
  n1(3 downto 3) &
  n1(2 downto 2) &
  n1(1 downto 1) &
  n1(0 downto 0);
process (clock_c) begin
  if rising_edge(clock_c) then
    if i5 = "1" then
      n4 <= "0000000000000000";
    elsif i4 = "1" then
      n4 <= i2;
    end if;
  end if;
end process;
n5 <= n4(15 downto 15) &
  n4(14 downto 14) &
  n4(13 downto 13) &
  n4(12 downto 12) &
  n4(11 downto 11) &
  n4(10 downto 10) &
  n4(9 downto 9) &
  n4(8 downto 8);
n6 <= n4(7 downto 7) &
  n4(6 downto 6) &
  n4(5 downto 5) &
  n4(4 downto 4) &
  n4(3 downto 3) &
  n4(2 downto 2) &
  n4(1 downto 1) &
  n4(0 downto 0);
process (clock_c) begin
  if rising_edge(clock_c) then
    if i5 = "1" then
      n7 <= "00000000";
    elsif i4 = "1" then
      n7 <= n2;
    end if;
  end if;
end process;
process (clock_c) begin
  if rising_edge(clock_c) then
    if i5 = "1" then
      n8 <= "00000000";
    elsif i4 = "1" then
      n8 <= n7;
    end if;
  end if;
end process;
process (clock_c) begin
  if rising_edge(clock_c) then
    if i5 = "1" then
      n9 <= "00000000";
    elsif i4 = "1" then
      n9 <= n3;
    end if;
  end if;
end process;
process (clock_c) begin
  if rising_edge(clock_c) then
    if i5 = "1" then
      n10 <= "00000000";
    elsif i4 = "1" then
      n10 <= n9;
    end if;
  end if;
end process;
process (clock_c) begin
  if rising_edge(clock_c) then 
    if i4 = "1" then
      case i3 is
        when "0000000" => n11 <= "0111111100000000";
        when "0000001" => n11 <= "0111111111111100";
        when "0000010" => n11 <= "0111111111111001";
        when "0000011" => n11 <= "0111111111110110";
        when "0000100" => n11 <= "0111111111110011";
        when "0000101" => n11 <= "0111111111110000";
        when "0000110" => n11 <= "0111111011101101";
        when "0000111" => n11 <= "0111111011101010";
        when "0001000" => n11 <= "0111110111100111";
        when "0001001" => n11 <= "0111110011100011";
        when "0001010" => n11 <= "0111110011100000";
        when "0001011" => n11 <= "0111101111011101";
        when "0001100" => n11 <= "0111101011011010";
        when "0001101" => n11 <= "0111100111010111";
        when "0001110" => n11 <= "0111100011010100";
        when "0001111" => n11 <= "0111011111010001";
        when "0010000" => n11 <= "0111011011001111";
        when "0010001" => n11 <= "0111010111001100";
        when "0010010" => n11 <= "0111001111001001";
        when "0010011" => n11 <= "0111001011000110";
        when "0010100" => n11 <= "0111000011000011";
        when "0010101" => n11 <= "0110111111000000";
        when "0010110" => n11 <= "0110110110111110";
        when "0010111" => n11 <= "0110110010111011";
        when "0011000" => n11 <= "0110101010111000";
        when "0011001" => n11 <= "0110100010110110";
        when "0011010" => n11 <= "0110011010110011";
        when "0011011" => n11 <= "0110010010110001";
        when "0011100" => n11 <= "0110001010101110";
        when "0011101" => n11 <= "0110000010101100";
        when "0011110" => n11 <= "0101111010101010";
        when "0011111" => n11 <= "0101110010100111";
        when "0100000" => n11 <= "0101101010100101";
        when "0100001" => n11 <= "0101100010100011";
        when "0100010" => n11 <= "0101010110100001";
        when "0100011" => n11 <= "0101001110011111";
        when "0100100" => n11 <= "0101000110011101";
        when "0100101" => n11 <= "0100111010011011";
        when "0100110" => n11 <= "0100110010011001";
        when "0100111" => n11 <= "0100100110010111";
        when "0101000" => n11 <= "0100011110010101";
        when "0101001" => n11 <= "0100010010010011";
        when "0101010" => n11 <= "0100000110010010";
        when "0101011" => n11 <= "0011111110010000";
        when "0101100" => n11 <= "0011110010001111";
        when "0101101" => n11 <= "0011100110001101";
        when "0101110" => n11 <= "0011011010001100";
        when "0101111" => n11 <= "0011001110001010";
        when "0110000" => n11 <= "0011000010001001";
        when "0110001" => n11 <= "0010111010001000";
        when "0110010" => n11 <= "0010101110000111";
        when "0110011" => n11 <= "0010100010000110";
        when "0110100" => n11 <= "0010010110000101";
        when "0110101" => n11 <= "0010001010000100";
        when "0110110" => n11 <= "0001111110000011";
        when "0110111" => n11 <= "0001110010000011";
        when "0111000" => n11 <= "0001100010000010";
        when "0111001" => n11 <= "0001010110000001";
        when "0111010" => n11 <= "0001001010000001";
        when "0111011" => n11 <= "0000111110000000";
        when "0111100" => n11 <= "0000110010000000";
        when "0111101" => n11 <= "0000100110000000";
        when "0111110" => n11 <= "0000011010000000";
        when "0111111" => n11 <= "0000001110000000";
        when "1000000" => n11 <= "0000000010000000";
        when "1000001" => n11 <= "1111110010000000";
        when "1000010" => n11 <= "1111100110000000";
        when "1000011" => n11 <= "1111011010000000";
        when "1000100" => n11 <= "1111001110000000";
        when "1000101" => n11 <= "1111000010000000";
        when "1000110" => n11 <= "1110110110000001";
        when "1000111" => n11 <= "1110101010000001";
        when "1001000" => n11 <= "1110011110000010";
        when "1001001" => n11 <= "1110001110000011";
        when "1001010" => n11 <= "1110000010000011";
        when "1001011" => n11 <= "1101110110000100";
        when "1001100" => n11 <= "1101101010000101";
        when "1001101" => n11 <= "1101011110000110";
        when "1001110" => n11 <= "1101010010000111";
        when "1001111" => n11 <= "1101000110001000";
        when "1010000" => n11 <= "1100111110001001";
        when "1010001" => n11 <= "1100110010001010";
        when "1010010" => n11 <= "1100100110001100";
        when "1010011" => n11 <= "1100011010001101";
        when "1010100" => n11 <= "1100001110001111";
        when "1010101" => n11 <= "1100000010010000";
        when "1010110" => n11 <= "1011111010010010";
        when "1010111" => n11 <= "1011101110010011";
        when "1011000" => n11 <= "1011100010010101";
        when "1011001" => n11 <= "1011011010010111";
        when "1011010" => n11 <= "1011001110011001";
        when "1011011" => n11 <= "1011000110011011";
        when "1011100" => n11 <= "1010111010011101";
        when "1011101" => n11 <= "1010110010011111";
        when "1011110" => n11 <= "1010101010100001";
        when "1011111" => n11 <= "1010011110100011";
        when "1100000" => n11 <= "1010010110100101";
        when "1100001" => n11 <= "1010001110100111";
        when "1100010" => n11 <= "1010000110101010";
        when "1100011" => n11 <= "1001111110101100";
        when "1100100" => n11 <= "1001110110101110";
        when "1100101" => n11 <= "1001101110110001";
        when "1100110" => n11 <= "1001100110110011";
        when "1100111" => n11 <= "1001011110110110";
        when "1101000" => n11 <= "1001010110111000";
        when "1101001" => n11 <= "1001001110111011";
        when "1101010" => n11 <= "1001001010111110";
        when "1101011" => n11 <= "1001000011000000";
        when "1101100" => n11 <= "1000111111000011";
        when "1101101" => n11 <= "1000110111000110";
        when "1101110" => n11 <= "1000110011001001";
        when "1101111" => n11 <= "1000101011001100";
        when "1110000" => n11 <= "1000100111001111";
        when "1110001" => n11 <= "1000100011010001";
        when "1110010" => n11 <= "1000011111010100";
        when "1110011" => n11 <= "1000011011010111";
        when "1110100" => n11 <= "1000010111011010";
        when "1110101" => n11 <= "1000010011011101";
        when "1110110" => n11 <= "1000001111100000";
        when "1110111" => n11 <= "1000001111100011";
        when "1111000" => n11 <= "1000001011100111";
        when "1111001" => n11 <= "1000000111101010";
        when "1111010" => n11 <= "1000000111101101";
        when "1111011" => n11 <= "1000000011110000";
        when "1111100" => n11 <= "1000000011110011";
        when "1111101" => n11 <= "1000000011110110";
        when "1111110" => n11 <= "1000000011111001";
        when "1111111" => n11 <= "1000000011111100";
        when others => n11 <= "XXXXXXXXXXXXXXXX";
      end case;
    end if;
  end if;
end process;
n12 <= n11(15 downto 15) &
  n11(14 downto 14) &
  n11(13 downto 13) &
  n11(12 downto 12) &
  n11(11 downto 11) &
  n11(10 downto 10) &
  n11(9 downto 9) &
  n11(8 downto 8);
n13 <= n11(7 downto 7) &
  n11(6 downto 6) &
  n11(5 downto 5) &
  n11(4 downto 4) &
  n11(3 downto 3) &
  n11(2 downto 2) &
  n11(1 downto 1) &
  n11(0 downto 0);
n14 <= unsigned(signed(n5) * signed(n12));
n15 <= n14(14 downto 14) &
  n14(13 downto 13) &
  n14(12 downto 12) &
  n14(11 downto 11) &
  n14(10 downto 10) &
  n14(9 downto 9) &
  n14(8 downto 8) &
  n14(7 downto 7);
process (clock_c) begin
  if rising_edge(clock_c) then
    if i5 = "1" then
      n16 <= "00000000";
    elsif i4 = "1" then
      n16 <= n15;
    end if;
  end if;
end process;
n17 <= unsigned(signed(n6) * signed(n13));
n18 <= n17(14 downto 14) &
  n17(13 downto 13) &
  n17(12 downto 12) &
  n17(11 downto 11) &
  n17(10 downto 10) &
  n17(9 downto 9) &
  n17(8 downto 8) &
  n17(7 downto 7);
process (clock_c) begin
  if rising_edge(clock_c) then
    if i5 = "1" then
      n19 <= "00000000";
    elsif i4 = "1" then
      n19 <= n18;
    end if;
  end if;
end process;
n20 <= n16 - n19;
process (clock_c) begin
  if rising_edge(clock_c) then
    if i5 = "1" then
      n21 <= "00000000";
    elsif i4 = "1" then
      n21 <= n20;
    end if;
  end if;
end process;
n22 <= unsigned(signed(n5) * signed(n13));
n23 <= n22(14 downto 14) &
  n22(13 downto 13) &
  n22(12 downto 12) &
  n22(11 downto 11) &
  n22(10 downto 10) &
  n22(9 downto 9) &
  n22(8 downto 8) &
  n22(7 downto 7);
process (clock_c) begin
  if rising_edge(clock_c) then
    if i5 = "1" then
      n24 <= "00000000";
    elsif i4 = "1" then
      n24 <= n23;
    end if;
  end if;
end process;
n25 <= unsigned(signed(n6) * signed(n12));
n26 <= n25(14 downto 14) &
  n25(13 downto 13) &
  n25(12 downto 12) &
  n25(11 downto 11) &
  n25(10 downto 10) &
  n25(9 downto 9) &
  n25(8 downto 8) &
  n25(7 downto 7);
process (clock_c) begin
  if rising_edge(clock_c) then
    if i5 = "1" then
      n27 <= "00000000";
    elsif i4 = "1" then
      n27 <= n26;
    end if;
  end if;
end process;
n28 <= n24 + n27;
process (clock_c) begin
  if rising_edge(clock_c) then
    if i5 = "1" then
      n29 <= "00000000";
    elsif i4 = "1" then
      n29 <= n28;
    end if;
  end if;
end process;
n30 <= n8 + n21;
n31 <= n10 + n29;
n32 <= n30 & n31;
process (clock_c) begin
  if rising_edge(clock_c) then
    if i5 = "1" then
      n33 <= "0000000000000000";
    elsif i4 = "1" then
      n33 <= n32;
    end if;
  end if;
end process;
n34 <= n8 - n21;
n35 <= n10 - n29;
n36 <= n34 & n35;
process (clock_c) begin
  if rising_edge(clock_c) then
    if i5 = "1" then
      n37 <= "0000000000000000";
    elsif i4 = "1" then
      n37 <= n36;
    end if;
  end if;
end process;
o2 <= n37;
o1 <= n33;
end architecture rtl;

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
entity cf_fft_2048_8_17 is
port (
clock_c : in std_logic;
i1 : in  unsigned(0 downto 0);
i2 : in  unsigned(15 downto 0);
i3 : in  unsigned(15 downto 0);
i4 : in  unsigned(0 downto 0);
i5 : in  unsigned(0 downto 0);
o1 : out unsigned(0 downto 0);
o2 : out unsigned(15 downto 0);
o3 : out unsigned(15 downto 0));
end entity cf_fft_2048_8_17;
architecture rtl of cf_fft_2048_8_17 is
signal n1 : unsigned(6 downto 0);
signal n2 : unsigned(31 downto 0);
signal n3 : unsigned(0 downto 0) := "0";
signal n4 : unsigned(0 downto 0) := "0";
signal n5 : unsigned(0 downto 0) := "0";
signal n6 : unsigned(0 downto 0) := "0";
signal n7 : unsigned(8 downto 0);
signal n8 : unsigned(8 downto 0) := "000000000";
signal n9 : unsigned(8 downto 0) := "000000000";
signal n10 : unsigned(8 downto 0) := "000000000";
signal n11 : unsigned(8 downto 0) := "000000000";
signal n12 : unsigned(0 downto 0);
signal n13 : unsigned(0 downto 0) := "0";
signal n14 : unsigned(0 downto 0) := "0";
signal n15 : unsigned(0 downto 0) := "0";
signal n16 : unsigned(0 downto 0) := "0";
signal n17 : unsigned(0 downto 0);
signal n18 : unsigned(1 downto 0);
signal n19 : unsigned(15 downto 0);
signal n20 : unsigned(15 downto 0);
signal n21 : unsigned(15 downto 0);
signal n22 : unsigned(15 downto 0);
signal n23 : unsigned(15 downto 0);
signal n24 : unsigned(15 downto 0);
signal s25_1 : unsigned(15 downto 0);
signal s25_2 : unsigned(15 downto 0);
signal s26_1 : unsigned(0 downto 0);
signal s27_1 : unsigned(9 downto 0);
signal s27_2 : unsigned(0 downto 0);
signal s28_1 : unsigned(31 downto 0);
signal s29_1 : unsigned(0 downto 0);
signal s29_2 : unsigned(0 downto 0);
signal s29_3 : unsigned(31 downto 0);
component cf_fft_2048_8_18 is
port (
clock_c : in std_logic;
i1 : in  unsigned(15 downto 0);
i2 : in  unsigned(15 downto 0);
i3 : in  unsigned(6 downto 0);
i4 : in  unsigned(0 downto 0);
i5 : in  unsigned(0 downto 0);
o1 : out unsigned(15 downto 0);
o2 : out unsigned(15 downto 0));
end component cf_fft_2048_8_18;
component cf_fft_2048_8_35 is
port (
clock_c : in std_logic;
i1 : in  unsigned(1 downto 0);
i2 : in  unsigned(0 downto 0);
i3 : in  unsigned(0 downto 0);
o1 : out unsigned(0 downto 0));
end component cf_fft_2048_8_35;
component cf_fft_2048_8_26 is
port (
clock_c : in std_logic;
i1 : in  unsigned(0 downto 0);
i2 : in  unsigned(0 downto 0);
i3 : in  unsigned(0 downto 0);
o1 : out unsigned(9 downto 0);
o2 : out unsigned(0 downto 0));
end component cf_fft_2048_8_26;
component cf_fft_2048_8_31 is
port (
clock_c : in std_logic;
i1 : in  unsigned(31 downto 0);
i2 : in  unsigned(0 downto 0);
i3 : in  unsigned(8 downto 0);
i4 : in  unsigned(0 downto 0);
i5 : in  unsigned(0 downto 0);
i6 : in  unsigned(0 downto 0);
o1 : out unsigned(31 downto 0));
end component cf_fft_2048_8_31;
component cf_fft_2048_8_30 is
port (
clock_c : in std_logic;
i1 : in  unsigned(31 downto 0);
i2 : in  unsigned(0 downto 0);
i3 : in  unsigned(8 downto 0);
i4 : in  unsigned(0 downto 0);
i5 : in  unsigned(0 downto 0);
i6 : in  unsigned(0 downto 0);
o1 : out unsigned(0 downto 0);
o2 : out unsigned(0 downto 0);
o3 : out unsigned(31 downto 0));
end component cf_fft_2048_8_30;
begin
n1 <= s27_1(9 downto 9) &
  s27_1(8 downto 8) &
  s27_1(7 downto 7) &
  s27_1(6 downto 6) &
  s27_1(5 downto 5) &
  s27_1(4 downto 4) &
  s27_1(3 downto 3);
n2 <= s25_1 & s25_2;
process (clock_c) begin
  if rising_edge(clock_c) then
    if i5 = "1" then
      n3 <= "0";
    elsif i4 = "1" then
      n3 <= s27_2;
    end if;
  end if;
end process;
process (clock_c) begin
  if rising_edge(clock_c) then
    if i5 = "1" then
      n4 <= "0";
    elsif i4 = "1" then
      n4 <= n3;
    end if;
  end if;
end process;
process (clock_c) begin
  if rising_edge(clock_c) then
    if i5 = "1" then
      n5 <= "0";
    elsif i4 = "1" then
      n5 <= n4;
    end if;
  end if;
end process;
process (clock_c) begin
  if rising_edge(clock_c) then
    if i5 = "1" then
      n6 <= "0";
    elsif i4 = "1" then
      n6 <= n5;
    end if;
  end if;
end process;
n7 <= s27_1(9 downto 9) &
  s27_1(8 downto 8) &
  s27_1(7 downto 7) &
  s27_1(6 downto 6) &
  s27_1(5 downto 5) &
  s27_1(4 downto 4) &
  s27_1(3 downto 3) &
  s27_1(2 downto 2) &
  s27_1(1 downto 1);
process (clock_c) begin
  if rising_edge(clock_c) then
    if i5 = "1" then
      n8 <= "000000000";
    elsif i4 = "1" then
      n8 <= n7;
    end if;
  end if;
end process;
process (clock_c) begin
  if rising_edge(clock_c) then
    if i5 = "1" then
      n9 <= "000000000";
    elsif i4 = "1" then
      n9 <= n8;
    end if;
  end if;
end process;
process (clock_c) begin
  if rising_edge(clock_c) then
    if i5 = "1" then
      n10 <= "000000000";
    elsif i4 = "1" then
      n10 <= n9;
    end if;
  end if;
end process;
process (clock_c) begin
  if rising_edge(clock_c) then
    if i5 = "1" then
      n11 <= "000000000";
    elsif i4 = "1" then
      n11 <= n10;
    end if;
  end if;
end process;
n12 <= s27_1(0 downto 0);
process (clock_c) begin
  if rising_edge(clock_c) then
    if i5 = "1" then
      n13 <= "0";
    elsif i4 = "1" then
      n13 <= n12;
    end if;
  end if;
end process;
process (clock_c) begin
  if rising_edge(clock_c) then
    if i5 = "1" then
      n14 <= "0";
    elsif i4 = "1" then
      n14 <= n13;
    end if;
  end if;
end process;
process (clock_c) begin
  if rising_edge(clock_c) then
    if i5 = "1" then
      n15 <= "0";
    elsif i4 = "1" then
      n15 <= n14;
    end if;
  end if;
end process;
process (clock_c) begin
  if rising_edge(clock_c) then
    if i5 = "1" then
      n16 <= "0";
    elsif i4 = "1" then
      n16 <= n15;
    end if;
  end if;
end process;
n17 <= not n16;
n18 <= s29_2 & s29_1;
n19 <= s29_3(31 downto 31) &
  s29_3(30 downto 30) &
  s29_3(29 downto 29) &
  s29_3(28 downto 28) &
  s29_3(27 downto 27) &
  s29_3(26 downto 26) &
  s29_3(25 downto 25) &
  s29_3(24 downto 24) &
  s29_3(23 downto 23) &
  s29_3(22 downto 22) &
  s29_3(21 downto 21) &
  s29_3(20 downto 20) &
  s29_3(19 downto 19) &
  s29_3(18 downto 18) &
  s29_3(17 downto 17) &
  s29_3(16 downto 16);
n20 <= s29_3(15 downto 15) &
  s29_3(14 downto 14) &
  s29_3(13 downto 13) &
  s29_3(12 downto 12) &
  s29_3(11 downto 11) &
  s29_3(10 downto 10) &
  s29_3(9 downto 9) &
  s29_3(8 downto 8) &
  s29_3(7 downto 7) &
  s29_3(6 downto 6) &
  s29_3(5 downto 5) &
  s29_3(4 downto 4) &
  s29_3(3 downto 3) &
  s29_3(2 downto 2) &
  s29_3(1 downto 1) &
  s29_3(0 downto 0);
n21 <= s28_1(31 downto 31) &
  s28_1(30 downto 30) &
  s28_1(29 downto 29) &
  s28_1(28 downto 28) &
  s28_1(27 downto 27) &
  s28_1(26 downto 26) &
  s28_1(25 downto 25) &
  s28_1(24 downto 24) &
  s28_1(23 downto 23) &
  s28_1(22 downto 22) &
  s28_1(21 downto 21) &
  s28_1(20 downto 20) &
  s28_1(19 downto 19) &
  s28_1(18 downto 18) &
  s28_1(17 downto 17) &
  s28_1(16 downto 16);
n22 <= s28_1(15 downto 15) &
  s28_1(14 downto 14) &
  s28_1(13 downto 13) &
  s28_1(12 downto 12) &
  s28_1(11 downto 11) &
  s28_1(10 downto 10) &
  s28_1(9 downto 9) &
  s28_1(8 downto 8) &
  s28_1(7 downto 7) &
  s28_1(6 downto 6) &
  s28_1(5 downto 5) &
  s28_1(4 downto 4) &
  s28_1(3 downto 3) &
  s28_1(2 downto 2) &
  s28_1(1 downto 1) &
  s28_1(0 downto 0);
n23 <= n20 when s26_1 = "1" else n19;
n24 <= n22 when s26_1 = "1" else n21;
s25 : cf_fft_2048_8_18 port map (clock_c, i2, i3, n1, i4, i5, s25_1, s25_2);
s26 : cf_fft_2048_8_35 port map (clock_c, n18, i4, i5, s26_1);
s27 : cf_fft_2048_8_26 port map (clock_c, i1, i4, i5, s27_1, s27_2);
s28 : cf_fft_2048_8_31 port map (clock_c, n2, n6, n11, n16, i4, i5, s28_1);
s29 : cf_fft_2048_8_30 port map (clock_c, n2, n6, n11, n17, i4, i5, s29_1, s29_2, s29_3);
o3 <= n24;
o2 <= n23;
o1 <= s29_1;
end architecture rtl;

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
entity cf_fft_2048_8_16 is
port (
clock_c : in std_logic;
i1 : in  unsigned(15 downto 0);
i2 : in  unsigned(15 downto 0);
i3 : in  unsigned(5 downto 0);
i4 : in  unsigned(0 downto 0);
i5 : in  unsigned(0 downto 0);
o1 : out unsigned(15 downto 0);
o2 : out unsigned(15 downto 0));
end entity cf_fft_2048_8_16;
architecture rtl of cf_fft_2048_8_16 is
signal n1 : unsigned(15 downto 0) := "0000000000000000";
signal n2 : unsigned(7 downto 0);
signal n3 : unsigned(7 downto 0);
signal n4 : unsigned(15 downto 0) := "0000000000000000";
signal n5 : unsigned(7 downto 0);
signal n6 : unsigned(7 downto 0);
signal n7 : unsigned(7 downto 0) := "00000000";
signal n8 : unsigned(7 downto 0) := "00000000";
signal n9 : unsigned(7 downto 0) := "00000000";
signal n10 : unsigned(7 downto 0) := "00000000";
signal n11 : unsigned(15 downto 0) := "0000000000000000";
signal n12 : unsigned(7 downto 0);
signal n13 : unsigned(7 downto 0);
signal n14 : unsigned(15 downto 0);
signal n15 : unsigned(7 downto 0);
signal n16 : unsigned(7 downto 0) := "00000000";
signal n17 : unsigned(15 downto 0);
signal n18 : unsigned(7 downto 0);
signal n19 : unsigned(7 downto 0) := "00000000";
signal n20 : unsigned(7 downto 0);
signal n21 : unsigned(7 downto 0) := "00000000";
signal n22 : unsigned(15 downto 0);
signal n23 : unsigned(7 downto 0);
signal n24 : unsigned(7 downto 0) := "00000000";
signal n25 : unsigned(15 downto 0);
signal n26 : unsigned(7 downto 0);
signal n27 : unsigned(7 downto 0) := "00000000";
signal n28 : unsigned(7 downto 0);
signal n29 : unsigned(7 downto 0) := "00000000";
signal n30 : unsigned(7 downto 0);
signal n31 : unsigned(7 downto 0);
signal n32 : unsigned(15 downto 0);
signal n33 : unsigned(15 downto 0) := "0000000000000000";
signal n34 : unsigned(7 downto 0);
signal n35 : unsigned(7 downto 0);
signal n36 : unsigned(15 downto 0);
signal n37 : unsigned(15 downto 0) := "0000000000000000";
begin
process (clock_c) begin
  if rising_edge(clock_c) then
    if i5 = "1" then
      n1 <= "0000000000000000";
    elsif i4 = "1" then
      n1 <= i1;
    end if;
  end if;
end process;
n2 <= n1(15 downto 15) &
  n1(14 downto 14) &
  n1(13 downto 13) &
  n1(12 downto 12) &
  n1(11 downto 11) &
  n1(10 downto 10) &
  n1(9 downto 9) &
  n1(8 downto 8);
n3 <= n1(7 downto 7) &
  n1(6 downto 6) &
  n1(5 downto 5) &
  n1(4 downto 4) &
  n1(3 downto 3) &
  n1(2 downto 2) &
  n1(1 downto 1) &
  n1(0 downto 0);
process (clock_c) begin
  if rising_edge(clock_c) then
    if i5 = "1" then
      n4 <= "0000000000000000";
    elsif i4 = "1" then
      n4 <= i2;
    end if;
  end if;
end process;
n5 <= n4(15 downto 15) &
  n4(14 downto 14) &
  n4(13 downto 13) &
  n4(12 downto 12) &
  n4(11 downto 11) &
  n4(10 downto 10) &
  n4(9 downto 9) &
  n4(8 downto 8);
n6 <= n4(7 downto 7) &
  n4(6 downto 6) &
  n4(5 downto 5) &
  n4(4 downto 4) &
  n4(3 downto 3) &
  n4(2 downto 2) &
  n4(1 downto 1) &
  n4(0 downto 0);
process (clock_c) begin
  if rising_edge(clock_c) then
    if i5 = "1" then
      n7 <= "00000000";
    elsif i4 = "1" then
      n7 <= n2;
    end if;
  end if;
end process;
process (clock_c) begin
  if rising_edge(clock_c) then
    if i5 = "1" then
      n8 <= "00000000";
    elsif i4 = "1" then
      n8 <= n7;
    end if;
  end if;
end process;
process (clock_c) begin
  if rising_edge(clock_c) then
    if i5 = "1" then
      n9 <= "00000000";
    elsif i4 = "1" then
      n9 <= n3;
    end if;
  end if;
end process;
process (clock_c) begin
  if rising_edge(clock_c) then
    if i5 = "1" then
      n10 <= "00000000";
    elsif i4 = "1" then
      n10 <= n9;
    end if;
  end if;
end process;
process (clock_c) begin
  if rising_edge(clock_c) then 
    if i4 = "1" then
      case i3 is
        when "000000" => n11 <= "0111111100000000";
        when "000001" => n11 <= "0111111111111001";
        when "000010" => n11 <= "0111111111110011";
        when "000011" => n11 <= "0111111011101101";
        when "000100" => n11 <= "0111110111100111";
        when "000101" => n11 <= "0111110011100000";
        when "000110" => n11 <= "0111101011011010";
        when "000111" => n11 <= "0111100011010100";
        when "001000" => n11 <= "0111011011001111";
        when "001001" => n11 <= "0111001111001001";
        when "001010" => n11 <= "0111000011000011";
        when "001011" => n11 <= "0110110110111110";
        when "001100" => n11 <= "0110101010111000";
        when "001101" => n11 <= "0110011010110011";
        when "001110" => n11 <= "0110001010101110";
        when "001111" => n11 <= "0101111010101010";
        when "010000" => n11 <= "0101101010100101";
        when "010001" => n11 <= "0101010110100001";
        when "010010" => n11 <= "0101000110011101";
        when "010011" => n11 <= "0100110010011001";
        when "010100" => n11 <= "0100011110010101";
        when "010101" => n11 <= "0100000110010010";
        when "010110" => n11 <= "0011110010001111";
        when "010111" => n11 <= "0011011010001100";
        when "011000" => n11 <= "0011000010001001";
        when "011001" => n11 <= "0010101110000111";
        when "011010" => n11 <= "0010010110000101";
        when "011011" => n11 <= "0001111110000011";
        when "011100" => n11 <= "0001100010000010";
        when "011101" => n11 <= "0001001010000001";
        when "011110" => n11 <= "0000110010000000";
        when "011111" => n11 <= "0000011010000000";
        when "100000" => n11 <= "0000000010000000";
        when "100001" => n11 <= "1111100110000000";
        when "100010" => n11 <= "1111001110000000";
        when "100011" => n11 <= "1110110110000001";
        when "100100" => n11 <= "1110011110000010";
        when "100101" => n11 <= "1110000010000011";
        when "100110" => n11 <= "1101101010000101";
        when "100111" => n11 <= "1101010010000111";
        when "101000" => n11 <= "1100111110001001";
        when "101001" => n11 <= "1100100110001100";
        when "101010" => n11 <= "1100001110001111";
        when "101011" => n11 <= "1011111010010010";
        when "101100" => n11 <= "1011100010010101";
        when "101101" => n11 <= "1011001110011001";
        when "101110" => n11 <= "1010111010011101";
        when "101111" => n11 <= "1010101010100001";
        when "110000" => n11 <= "1010010110100101";
        when "110001" => n11 <= "1010000110101010";
        when "110010" => n11 <= "1001110110101110";
        when "110011" => n11 <= "1001100110110011";
        when "110100" => n11 <= "1001010110111000";
        when "110101" => n11 <= "1001001010111110";
        when "110110" => n11 <= "1000111111000011";
        when "110111" => n11 <= "1000110011001001";
        when "111000" => n11 <= "1000100111001111";
        when "111001" => n11 <= "1000011111010100";
        when "111010" => n11 <= "1000010111011010";
        when "111011" => n11 <= "1000001111100000";
        when "111100" => n11 <= "1000001011100111";
        when "111101" => n11 <= "1000000111101101";
        when "111110" => n11 <= "1000000011110011";
        when "111111" => n11 <= "1000000011111001";
        when others => n11 <= "XXXXXXXXXXXXXXXX";
      end case;
    end if;
  end if;
end process;
n12 <= n11(15 downto 15) &
  n11(14 downto 14) &
  n11(13 downto 13) &
  n11(12 downto 12) &
  n11(11 downto 11) &
  n11(10 downto 10) &
  n11(9 downto 9) &
  n11(8 downto 8);
n13 <= n11(7 downto 7) &
  n11(6 downto 6) &
  n11(5 downto 5) &
  n11(4 downto 4) &
  n11(3 downto 3) &
  n11(2 downto 2) &
  n11(1 downto 1) &
  n11(0 downto 0);
n14 <= unsigned(signed(n5) * signed(n12));
n15 <= n14(14 downto 14) &
  n14(13 downto 13) &
  n14(12 downto 12) &
  n14(11 downto 11) &
  n14(10 downto 10) &
  n14(9 downto 9) &
  n14(8 downto 8) &
  n14(7 downto 7);
process (clock_c) begin
  if rising_edge(clock_c) then
    if i5 = "1" then
      n16 <= "00000000";
    elsif i4 = "1" then
      n16 <= n15;
    end if;
  end if;
end process;
n17 <= unsigned(signed(n6) * signed(n13));
n18 <= n17(14 downto 14) &
  n17(13 downto 13) &
  n17(12 downto 12) &
  n17(11 downto 11) &
  n17(10 downto 10) &
  n17(9 downto 9) &
  n17(8 downto 8) &
  n17(7 downto 7);
process (clock_c) begin
  if rising_edge(clock_c) then
    if i5 = "1" then
      n19 <= "00000000";
    elsif i4 = "1" then
      n19 <= n18;
    end if;
  end if;
end process;
n20 <= n16 - n19;
process (clock_c) begin
  if rising_edge(clock_c) then
    if i5 = "1" then
      n21 <= "00000000";
    elsif i4 = "1" then
      n21 <= n20;
    end if;
  end if;
end process;
n22 <= unsigned(signed(n5) * signed(n13));
n23 <= n22(14 downto 14) &
  n22(13 downto 13) &
  n22(12 downto 12) &
  n22(11 downto 11) &
  n22(10 downto 10) &
  n22(9 downto 9) &
  n22(8 downto 8) &
  n22(7 downto 7);
process (clock_c) begin
  if rising_edge(clock_c) then
    if i5 = "1" then
      n24 <= "00000000";
    elsif i4 = "1" then
      n24 <= n23;
    end if;
  end if;
end process;
n25 <= unsigned(signed(n6) * signed(n12));
n26 <= n25(14 downto 14) &
  n25(13 downto 13) &
  n25(12 downto 12) &
  n25(11 downto 11) &
  n25(10 downto 10) &
  n25(9 downto 9) &
  n25(8 downto 8) &
  n25(7 downto 7);
process (clock_c) begin
  if rising_edge(clock_c) then
    if i5 = "1" then
      n27 <= "00000000";
    elsif i4 = "1" then
      n27 <= n26;
    end if;
  end if;
end process;
n28 <= n24 + n27;
process (clock_c) begin
  if rising_edge(clock_c) then
    if i5 = "1" then
      n29 <= "00000000";
    elsif i4 = "1" then
      n29 <= n28;
    end if;
  end if;
end process;
n30 <= n8 + n21;
n31 <= n10 + n29;
n32 <= n30 & n31;
process (clock_c) begin
  if rising_edge(clock_c) then
    if i5 = "1" then
      n33 <= "0000000000000000";
    elsif i4 = "1" then
      n33 <= n32;
    end if;
  end if;
end process;
n34 <= n8 - n21;
n35 <= n10 - n29;
n36 <= n34 & n35;
process (clock_c) begin
  if rising_edge(clock_c) then
    if i5 = "1" then
      n37 <= "0000000000000000";
    elsif i4 = "1" then
      n37 <= n36;
    end if;
  end if;
end process;
o2 <= n37;
o1 <= n33;
end architecture rtl;

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
entity cf_fft_2048_8_15 is
port (
clock_c : in std_logic;
i1 : in  unsigned(0 downto 0);
i2 : in  unsigned(15 downto 0);
i3 : in  unsigned(15 downto 0);
i4 : in  unsigned(0 downto 0);
i5 : in  unsigned(0 downto 0);
o1 : out unsigned(0 downto 0);
o2 : out unsigned(15 downto 0);
o3 : out unsigned(15 downto 0));
end entity cf_fft_2048_8_15;
architecture rtl of cf_fft_2048_8_15 is
signal n1 : unsigned(5 downto 0);
signal n2 : unsigned(31 downto 0);
signal n3 : unsigned(0 downto 0) := "0";
signal n4 : unsigned(0 downto 0) := "0";
signal n5 : unsigned(0 downto 0) := "0";
signal n6 : unsigned(0 downto 0) := "0";
signal n7 : unsigned(8 downto 0);
signal n8 : unsigned(8 downto 0) := "000000000";
signal n9 : unsigned(8 downto 0) := "000000000";
signal n10 : unsigned(8 downto 0) := "000000000";
signal n11 : unsigned(8 downto 0) := "000000000";
signal n12 : unsigned(0 downto 0);
signal n13 : unsigned(0 downto 0) := "0";
signal n14 : unsigned(0 downto 0) := "0";
signal n15 : unsigned(0 downto 0) := "0";
signal n16 : unsigned(0 downto 0) := "0";
signal n17 : unsigned(0 downto 0);
signal n18 : unsigned(1 downto 0);
signal n19 : unsigned(15 downto 0);
signal n20 : unsigned(15 downto 0);
signal n21 : unsigned(15 downto 0);
signal n22 : unsigned(15 downto 0);
signal n23 : unsigned(15 downto 0);
signal n24 : unsigned(15 downto 0);
signal s25_1 : unsigned(0 downto 0);
signal s26_1 : unsigned(15 downto 0);
signal s26_2 : unsigned(15 downto 0);
signal s27_1 : unsigned(9 downto 0);
signal s27_2 : unsigned(0 downto 0);
signal s28_1 : unsigned(0 downto 0);
signal s28_2 : unsigned(0 downto 0);
signal s28_3 : unsigned(31 downto 0);
signal s29_1 : unsigned(31 downto 0);
component cf_fft_2048_8_35 is
port (
clock_c : in std_logic;
i1 : in  unsigned(1 downto 0);
i2 : in  unsigned(0 downto 0);
i3 : in  unsigned(0 downto 0);
o1 : out unsigned(0 downto 0));
end component cf_fft_2048_8_35;
component cf_fft_2048_8_16 is
port (
clock_c : in std_logic;
i1 : in  unsigned(15 downto 0);
i2 : in  unsigned(15 downto 0);
i3 : in  unsigned(5 downto 0);
i4 : in  unsigned(0 downto 0);
i5 : in  unsigned(0 downto 0);
o1 : out unsigned(15 downto 0);
o2 : out unsigned(15 downto 0));
end component cf_fft_2048_8_16;
component cf_fft_2048_8_26 is
port (
clock_c : in std_logic;
i1 : in  unsigned(0 downto 0);
i2 : in  unsigned(0 downto 0);
i3 : in  unsigned(0 downto 0);
o1 : out unsigned(9 downto 0);
o2 : out unsigned(0 downto 0));
end component cf_fft_2048_8_26;
component cf_fft_2048_8_30 is
port (
clock_c : in std_logic;
i1 : in  unsigned(31 downto 0);
i2 : in  unsigned(0 downto 0);
i3 : in  unsigned(8 downto 0);
i4 : in  unsigned(0 downto 0);
i5 : in  unsigned(0 downto 0);
i6 : in  unsigned(0 downto 0);
o1 : out unsigned(0 downto 0);
o2 : out unsigned(0 downto 0);
o3 : out unsigned(31 downto 0));
end component cf_fft_2048_8_30;
component cf_fft_2048_8_31 is
port (
clock_c : in std_logic;
i1 : in  unsigned(31 downto 0);
i2 : in  unsigned(0 downto 0);
i3 : in  unsigned(8 downto 0);
i4 : in  unsigned(0 downto 0);
i5 : in  unsigned(0 downto 0);
i6 : in  unsigned(0 downto 0);
o1 : out unsigned(31 downto 0));
end component cf_fft_2048_8_31;
begin
n1 <= s27_1(9 downto 9) &
  s27_1(8 downto 8) &
  s27_1(7 downto 7) &
  s27_1(6 downto 6) &
  s27_1(5 downto 5) &
  s27_1(4 downto 4);
n2 <= s26_1 & s26_2;
process (clock_c) begin
  if rising_edge(clock_c) then
    if i5 = "1" then
      n3 <= "0";
    elsif i4 = "1" then
      n3 <= s27_2;
    end if;
  end if;
end process;
process (clock_c) begin
  if rising_edge(clock_c) then
    if i5 = "1" then
      n4 <= "0";
    elsif i4 = "1" then
      n4 <= n3;
    end if;
  end if;
end process;
process (clock_c) begin
  if rising_edge(clock_c) then
    if i5 = "1" then
      n5 <= "0";
    elsif i4 = "1" then
      n5 <= n4;
    end if;
  end if;
end process;
process (clock_c) begin
  if rising_edge(clock_c) then
    if i5 = "1" then
      n6 <= "0";
    elsif i4 = "1" then
      n6 <= n5;
    end if;
  end if;
end process;
n7 <= s27_1(9 downto 9) &
  s27_1(8 downto 8) &
  s27_1(7 downto 7) &
  s27_1(6 downto 6) &
  s27_1(5 downto 5) &
  s27_1(4 downto 4) &
  s27_1(3 downto 3) &
  s27_1(2 downto 2) &
  s27_1(1 downto 1);
process (clock_c) begin
  if rising_edge(clock_c) then
    if i5 = "1" then
      n8 <= "000000000";
    elsif i4 = "1" then
      n8 <= n7;
    end if;
  end if;
end process;
process (clock_c) begin
  if rising_edge(clock_c) then
    if i5 = "1" then
      n9 <= "000000000";
    elsif i4 = "1" then
      n9 <= n8;
    end if;
  end if;
end process;
process (clock_c) begin
  if rising_edge(clock_c) then
    if i5 = "1" then
      n10 <= "000000000";
    elsif i4 = "1" then
      n10 <= n9;
    end if;
  end if;
end process;
process (clock_c) begin
  if rising_edge(clock_c) then
    if i5 = "1" then
      n11 <= "000000000";
    elsif i4 = "1" then
      n11 <= n10;
    end if;
  end if;
end process;
n12 <= s27_1(0 downto 0);
process (clock_c) begin
  if rising_edge(clock_c) then
    if i5 = "1" then
      n13 <= "0";
    elsif i4 = "1" then
      n13 <= n12;
    end if;
  end if;
end process;
process (clock_c) begin
  if rising_edge(clock_c) then
    if i5 = "1" then
      n14 <= "0";
    elsif i4 = "1" then
      n14 <= n13;
    end if;
  end if;
end process;
process (clock_c) begin
  if rising_edge(clock_c) then
    if i5 = "1" then
      n15 <= "0";
    elsif i4 = "1" then
      n15 <= n14;
    end if;
  end if;
end process;
process (clock_c) begin
  if rising_edge(clock_c) then
    if i5 = "1" then
      n16 <= "0";
    elsif i4 = "1" then
      n16 <= n15;
    end if;
  end if;
end process;
n17 <= not n16;
n18 <= s28_2 & s28_1;
n19 <= s28_3(31 downto 31) &
  s28_3(30 downto 30) &
  s28_3(29 downto 29) &
  s28_3(28 downto 28) &
  s28_3(27 downto 27) &
  s28_3(26 downto 26) &
  s28_3(25 downto 25) &
  s28_3(24 downto 24) &
  s28_3(23 downto 23) &
  s28_3(22 downto 22) &
  s28_3(21 downto 21) &
  s28_3(20 downto 20) &
  s28_3(19 downto 19) &
  s28_3(18 downto 18) &
  s28_3(17 downto 17) &
  s28_3(16 downto 16);
n20 <= s28_3(15 downto 15) &
  s28_3(14 downto 14) &
  s28_3(13 downto 13) &
  s28_3(12 downto 12) &
  s28_3(11 downto 11) &
  s28_3(10 downto 10) &
  s28_3(9 downto 9) &
  s28_3(8 downto 8) &
  s28_3(7 downto 7) &
  s28_3(6 downto 6) &
  s28_3(5 downto 5) &
  s28_3(4 downto 4) &
  s28_3(3 downto 3) &
  s28_3(2 downto 2) &
  s28_3(1 downto 1) &
  s28_3(0 downto 0);
n21 <= s29_1(31 downto 31) &
  s29_1(30 downto 30) &
  s29_1(29 downto 29) &
  s29_1(28 downto 28) &
  s29_1(27 downto 27) &
  s29_1(26 downto 26) &
  s29_1(25 downto 25) &
  s29_1(24 downto 24) &
  s29_1(23 downto 23) &
  s29_1(22 downto 22) &
  s29_1(21 downto 21) &
  s29_1(20 downto 20) &
  s29_1(19 downto 19) &
  s29_1(18 downto 18) &
  s29_1(17 downto 17) &
  s29_1(16 downto 16);
n22 <= s29_1(15 downto 15) &
  s29_1(14 downto 14) &
  s29_1(13 downto 13) &
  s29_1(12 downto 12) &
  s29_1(11 downto 11) &
  s29_1(10 downto 10) &
  s29_1(9 downto 9) &
  s29_1(8 downto 8) &
  s29_1(7 downto 7) &
  s29_1(6 downto 6) &
  s29_1(5 downto 5) &
  s29_1(4 downto 4) &
  s29_1(3 downto 3) &
  s29_1(2 downto 2) &
  s29_1(1 downto 1) &
  s29_1(0 downto 0);
n23 <= n20 when s25_1 = "1" else n19;
n24 <= n22 when s25_1 = "1" else n21;
s25 : cf_fft_2048_8_35 port map (clock_c, n18, i4, i5, s25_1);
s26 : cf_fft_2048_8_16 port map (clock_c, i2, i3, n1, i4, i5, s26_1, s26_2);
s27 : cf_fft_2048_8_26 port map (clock_c, i1, i4, i5, s27_1, s27_2);
s28 : cf_fft_2048_8_30 port map (clock_c, n2, n6, n11, n17, i4, i5, s28_1, s28_2, s28_3);
s29 : cf_fft_2048_8_31 port map (clock_c, n2, n6, n11, n16, i4, i5, s29_1);
o3 <= n24;
o2 <= n23;
o1 <= s28_1;
end architecture rtl;

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
entity cf_fft_2048_8_14 is
port (
clock_c : in std_logic;
i1 : in  unsigned(15 downto 0);
i2 : in  unsigned(15 downto 0);
i3 : in  unsigned(4 downto 0);
i4 : in  unsigned(0 downto 0);
i5 : in  unsigned(0 downto 0);
o1 : out unsigned(15 downto 0);
o2 : out unsigned(15 downto 0));
end entity cf_fft_2048_8_14;
architecture rtl of cf_fft_2048_8_14 is
signal n1 : unsigned(15 downto 0) := "0000000000000000";
signal n2 : unsigned(7 downto 0);
signal n3 : unsigned(7 downto 0);
signal n4 : unsigned(15 downto 0) := "0000000000000000";
signal n5 : unsigned(7 downto 0);
signal n6 : unsigned(7 downto 0);
signal n7 : unsigned(7 downto 0) := "00000000";
signal n8 : unsigned(7 downto 0) := "00000000";
signal n9 : unsigned(7 downto 0) := "00000000";
signal n10 : unsigned(7 downto 0) := "00000000";
signal n11 : unsigned(15 downto 0) := "0000000000000000";
signal n12 : unsigned(7 downto 0);
signal n13 : unsigned(7 downto 0);
signal n14 : unsigned(15 downto 0);
signal n15 : unsigned(7 downto 0);
signal n16 : unsigned(7 downto 0) := "00000000";
signal n17 : unsigned(15 downto 0);
signal n18 : unsigned(7 downto 0);
signal n19 : unsigned(7 downto 0) := "00000000";
signal n20 : unsigned(7 downto 0);
signal n21 : unsigned(7 downto 0) := "00000000";
signal n22 : unsigned(15 downto 0);
signal n23 : unsigned(7 downto 0);
signal n24 : unsigned(7 downto 0) := "00000000";
signal n25 : unsigned(15 downto 0);
signal n26 : unsigned(7 downto 0);
signal n27 : unsigned(7 downto 0) := "00000000";
signal n28 : unsigned(7 downto 0);
signal n29 : unsigned(7 downto 0) := "00000000";
signal n30 : unsigned(7 downto 0);
signal n31 : unsigned(7 downto 0);
signal n32 : unsigned(15 downto 0);
signal n33 : unsigned(15 downto 0) := "0000000000000000";
signal n34 : unsigned(7 downto 0);
signal n35 : unsigned(7 downto 0);
signal n36 : unsigned(15 downto 0);
signal n37 : unsigned(15 downto 0) := "0000000000000000";
begin
process (clock_c) begin
  if rising_edge(clock_c) then
    if i5 = "1" then
      n1 <= "0000000000000000";
    elsif i4 = "1" then
      n1 <= i1;
    end if;
  end if;
end process;
n2 <= n1(15 downto 15) &
  n1(14 downto 14) &
  n1(13 downto 13) &
  n1(12 downto 12) &
  n1(11 downto 11) &
  n1(10 downto 10) &
  n1(9 downto 9) &
  n1(8 downto 8);
n3 <= n1(7 downto 7) &
  n1(6 downto 6) &
  n1(5 downto 5) &
  n1(4 downto 4) &
  n1(3 downto 3) &
  n1(2 downto 2) &
  n1(1 downto 1) &
  n1(0 downto 0);
process (clock_c) begin
  if rising_edge(clock_c) then
    if i5 = "1" then
      n4 <= "0000000000000000";
    elsif i4 = "1" then
      n4 <= i2;
    end if;
  end if;
end process;
n5 <= n4(15 downto 15) &
  n4(14 downto 14) &
  n4(13 downto 13) &
  n4(12 downto 12) &
  n4(11 downto 11) &
  n4(10 downto 10) &
  n4(9 downto 9) &
  n4(8 downto 8);
n6 <= n4(7 downto 7) &
  n4(6 downto 6) &
  n4(5 downto 5) &
  n4(4 downto 4) &
  n4(3 downto 3) &
  n4(2 downto 2) &
  n4(1 downto 1) &
  n4(0 downto 0);
process (clock_c) begin
  if rising_edge(clock_c) then
    if i5 = "1" then
      n7 <= "00000000";
    elsif i4 = "1" then
      n7 <= n2;
    end if;
  end if;
end process;
process (clock_c) begin
  if rising_edge(clock_c) then
    if i5 = "1" then
      n8 <= "00000000";
    elsif i4 = "1" then
      n8 <= n7;
    end if;
  end if;
end process;
process (clock_c) begin
  if rising_edge(clock_c) then
    if i5 = "1" then
      n9 <= "00000000";
    elsif i4 = "1" then
      n9 <= n3;
    end if;
  end if;
end process;
process (clock_c) begin
  if rising_edge(clock_c) then
    if i5 = "1" then
      n10 <= "00000000";
    elsif i4 = "1" then
      n10 <= n9;
    end if;
  end if;
end process;
process (clock_c) begin
  if rising_edge(clock_c) then 
    if i4 = "1" then
      case i3 is
        when "00000" => n11 <= "0111111100000000";
        when "00001" => n11 <= "0111111111110011";
        when "00010" => n11 <= "0111110111100111";
        when "00011" => n11 <= "0111101011011010";
        when "00100" => n11 <= "0111011011001111";
        when "00101" => n11 <= "0111000011000011";
        when "00110" => n11 <= "0110101010111000";
        when "00111" => n11 <= "0110001010101110";
        when "01000" => n11 <= "0101101010100101";
        when "01001" => n11 <= "0101000110011101";
        when "01010" => n11 <= "0100011110010101";
        when "01011" => n11 <= "0011110010001111";
        when "01100" => n11 <= "0011000010001001";
        when "01101" => n11 <= "0010010110000101";
        when "01110" => n11 <= "0001100010000010";
        when "01111" => n11 <= "0000110010000000";
        when "10000" => n11 <= "0000000010000000";
        when "10001" => n11 <= "1111001110000000";
        when "10010" => n11 <= "1110011110000010";
        when "10011" => n11 <= "1101101010000101";
        when "10100" => n11 <= "1100111110001001";
        when "10101" => n11 <= "1100001110001111";
        when "10110" => n11 <= "1011100010010101";
        when "10111" => n11 <= "1010111010011101";
        when "11000" => n11 <= "1010010110100101";
        when "11001" => n11 <= "1001110110101110";
        when "11010" => n11 <= "1001010110111000";
        when "11011" => n11 <= "1000111111000011";
        when "11100" => n11 <= "1000100111001111";
        when "11101" => n11 <= "1000010111011010";
        when "11110" => n11 <= "1000001011100111";
        when "11111" => n11 <= "1000000011110011";
        when others => n11 <= "XXXXXXXXXXXXXXXX";
      end case;
    end if;
  end if;
end process;
n12 <= n11(15 downto 15) &
  n11(14 downto 14) &
  n11(13 downto 13) &
  n11(12 downto 12) &
  n11(11 downto 11) &
  n11(10 downto 10) &
  n11(9 downto 9) &
  n11(8 downto 8);
n13 <= n11(7 downto 7) &
  n11(6 downto 6) &
  n11(5 downto 5) &
  n11(4 downto 4) &
  n11(3 downto 3) &
  n11(2 downto 2) &
  n11(1 downto 1) &
  n11(0 downto 0);
n14 <= unsigned(signed(n5) * signed(n12));
n15 <= n14(14 downto 14) &
  n14(13 downto 13) &
  n14(12 downto 12) &
  n14(11 downto 11) &
  n14(10 downto 10) &
  n14(9 downto 9) &
  n14(8 downto 8) &
  n14(7 downto 7);
process (clock_c) begin
  if rising_edge(clock_c) then
    if i5 = "1" then
      n16 <= "00000000";
    elsif i4 = "1" then
      n16 <= n15;
    end if;
  end if;
end process;
n17 <= unsigned(signed(n6) * signed(n13));
n18 <= n17(14 downto 14) &
  n17(13 downto 13) &
  n17(12 downto 12) &
  n17(11 downto 11) &
  n17(10 downto 10) &
  n17(9 downto 9) &
  n17(8 downto 8) &
  n17(7 downto 7);
process (clock_c) begin
  if rising_edge(clock_c) then
    if i5 = "1" then
      n19 <= "00000000";
    elsif i4 = "1" then
      n19 <= n18;
    end if;
  end if;
end process;
n20 <= n16 - n19;
process (clock_c) begin
  if rising_edge(clock_c) then
    if i5 = "1" then
      n21 <= "00000000";
    elsif i4 = "1" then
      n21 <= n20;
    end if;
  end if;
end process;
n22 <= unsigned(signed(n5) * signed(n13));
n23 <= n22(14 downto 14) &
  n22(13 downto 13) &
  n22(12 downto 12) &
  n22(11 downto 11) &
  n22(10 downto 10) &
  n22(9 downto 9) &
  n22(8 downto 8) &
  n22(7 downto 7);
process (clock_c) begin
  if rising_edge(clock_c) then
    if i5 = "1" then
      n24 <= "00000000";
    elsif i4 = "1" then
      n24 <= n23;
    end if;
  end if;
end process;
n25 <= unsigned(signed(n6) * signed(n12));
n26 <= n25(14 downto 14) &
  n25(13 downto 13) &
  n25(12 downto 12) &
  n25(11 downto 11) &
  n25(10 downto 10) &
  n25(9 downto 9) &
  n25(8 downto 8) &
  n25(7 downto 7);
process (clock_c) begin
  if rising_edge(clock_c) then
    if i5 = "1" then
      n27 <= "00000000";
    elsif i4 = "1" then
      n27 <= n26;
    end if;
  end if;
end process;
n28 <= n24 + n27;
process (clock_c) begin
  if rising_edge(clock_c) then
    if i5 = "1" then
      n29 <= "00000000";
    elsif i4 = "1" then
      n29 <= n28;
    end if;
  end if;
end process;
n30 <= n8 + n21;
n31 <= n10 + n29;
n32 <= n30 & n31;
process (clock_c) begin
  if rising_edge(clock_c) then
    if i5 = "1" then
      n33 <= "0000000000000000";
    elsif i4 = "1" then
      n33 <= n32;
    end if;
  end if;
end process;
n34 <= n8 - n21;
n35 <= n10 - n29;
n36 <= n34 & n35;
process (clock_c) begin
  if rising_edge(clock_c) then
    if i5 = "1" then
      n37 <= "0000000000000000";
    elsif i4 = "1" then
      n37 <= n36;
    end if;
  end if;
end process;
o2 <= n37;
o1 <= n33;
end architecture rtl;

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
entity cf_fft_2048_8_13 is
port (
clock_c : in std_logic;
i1 : in  unsigned(0 downto 0);
i2 : in  unsigned(15 downto 0);
i3 : in  unsigned(15 downto 0);
i4 : in  unsigned(0 downto 0);
i5 : in  unsigned(0 downto 0);
o1 : out unsigned(0 downto 0);
o2 : out unsigned(15 downto 0);
o3 : out unsigned(15 downto 0));
end entity cf_fft_2048_8_13;
architecture rtl of cf_fft_2048_8_13 is
signal n1 : unsigned(4 downto 0);
signal n2 : unsigned(31 downto 0);
signal n3 : unsigned(0 downto 0) := "0";
signal n4 : unsigned(0 downto 0) := "0";
signal n5 : unsigned(0 downto 0) := "0";
signal n6 : unsigned(0 downto 0) := "0";
signal n7 : unsigned(8 downto 0);
signal n8 : unsigned(8 downto 0) := "000000000";
signal n9 : unsigned(8 downto 0) := "000000000";
signal n10 : unsigned(8 downto 0) := "000000000";
signal n11 : unsigned(8 downto 0) := "000000000";
signal n12 : unsigned(0 downto 0);
signal n13 : unsigned(0 downto 0) := "0";
signal n14 : unsigned(0 downto 0) := "0";
signal n15 : unsigned(0 downto 0) := "0";
signal n16 : unsigned(0 downto 0) := "0";
signal n17 : unsigned(0 downto 0);
signal n18 : unsigned(1 downto 0);
signal n19 : unsigned(15 downto 0);
signal n20 : unsigned(15 downto 0);
signal n21 : unsigned(15 downto 0);
signal n22 : unsigned(15 downto 0);
signal n23 : unsigned(15 downto 0);
signal n24 : unsigned(15 downto 0);
signal s25_1 : unsigned(0 downto 0);
signal s26_1 : unsigned(15 downto 0);
signal s26_2 : unsigned(15 downto 0);
signal s27_1 : unsigned(9 downto 0);
signal s27_2 : unsigned(0 downto 0);
signal s28_1 : unsigned(0 downto 0);
signal s28_2 : unsigned(0 downto 0);
signal s28_3 : unsigned(31 downto 0);
signal s29_1 : unsigned(31 downto 0);
component cf_fft_2048_8_35 is
port (
clock_c : in std_logic;
i1 : in  unsigned(1 downto 0);
i2 : in  unsigned(0 downto 0);
i3 : in  unsigned(0 downto 0);
o1 : out unsigned(0 downto 0));
end component cf_fft_2048_8_35;
component cf_fft_2048_8_14 is
port (
clock_c : in std_logic;
i1 : in  unsigned(15 downto 0);
i2 : in  unsigned(15 downto 0);
i3 : in  unsigned(4 downto 0);
i4 : in  unsigned(0 downto 0);
i5 : in  unsigned(0 downto 0);
o1 : out unsigned(15 downto 0);
o2 : out unsigned(15 downto 0));
end component cf_fft_2048_8_14;
component cf_fft_2048_8_26 is
port (
clock_c : in std_logic;
i1 : in  unsigned(0 downto 0);
i2 : in  unsigned(0 downto 0);
i3 : in  unsigned(0 downto 0);
o1 : out unsigned(9 downto 0);
o2 : out unsigned(0 downto 0));
end component cf_fft_2048_8_26;
component cf_fft_2048_8_30 is
port (
clock_c : in std_logic;
i1 : in  unsigned(31 downto 0);
i2 : in  unsigned(0 downto 0);
i3 : in  unsigned(8 downto 0);
i4 : in  unsigned(0 downto 0);
i5 : in  unsigned(0 downto 0);
i6 : in  unsigned(0 downto 0);
o1 : out unsigned(0 downto 0);
o2 : out unsigned(0 downto 0);
o3 : out unsigned(31 downto 0));
end component cf_fft_2048_8_30;
component cf_fft_2048_8_31 is
port (
clock_c : in std_logic;
i1 : in  unsigned(31 downto 0);
i2 : in  unsigned(0 downto 0);
i3 : in  unsigned(8 downto 0);
i4 : in  unsigned(0 downto 0);
i5 : in  unsigned(0 downto 0);
i6 : in  unsigned(0 downto 0);
o1 : out unsigned(31 downto 0));
end component cf_fft_2048_8_31;
begin
n1 <= s27_1(9 downto 9) &
  s27_1(8 downto 8) &
  s27_1(7 downto 7) &
  s27_1(6 downto 6) &
  s27_1(5 downto 5);
n2 <= s26_1 & s26_2;
process (clock_c) begin
  if rising_edge(clock_c) then
    if i5 = "1" then
      n3 <= "0";
    elsif i4 = "1" then
      n3 <= s27_2;
    end if;
  end if;
end process;
process (clock_c) begin
  if rising_edge(clock_c) then
    if i5 = "1" then
      n4 <= "0";
    elsif i4 = "1" then
      n4 <= n3;
    end if;
  end if;
end process;
process (clock_c) begin
  if rising_edge(clock_c) then
    if i5 = "1" then
      n5 <= "0";
    elsif i4 = "1" then
      n5 <= n4;
    end if;
  end if;
end process;
process (clock_c) begin
  if rising_edge(clock_c) then
    if i5 = "1" then
      n6 <= "0";
    elsif i4 = "1" then
      n6 <= n5;
    end if;
  end if;
end process;
n7 <= s27_1(9 downto 9) &
  s27_1(8 downto 8) &
  s27_1(7 downto 7) &
  s27_1(6 downto 6) &
  s27_1(5 downto 5) &
  s27_1(4 downto 4) &
  s27_1(3 downto 3) &
  s27_1(2 downto 2) &
  s27_1(1 downto 1);
process (clock_c) begin
  if rising_edge(clock_c) then
    if i5 = "1" then
      n8 <= "000000000";
    elsif i4 = "1" then
      n8 <= n7;
    end if;
  end if;
end process;
process (clock_c) begin
  if rising_edge(clock_c) then
    if i5 = "1" then
      n9 <= "000000000";
    elsif i4 = "1" then
      n9 <= n8;
    end if;
  end if;
end process;
process (clock_c) begin
  if rising_edge(clock_c) then
    if i5 = "1" then
      n10 <= "000000000";
    elsif i4 = "1" then
      n10 <= n9;
    end if;
  end if;
end process;
process (clock_c) begin
  if rising_edge(clock_c) then
    if i5 = "1" then
      n11 <= "000000000";
    elsif i4 = "1" then
      n11 <= n10;
    end if;
  end if;
end process;
n12 <= s27_1(0 downto 0);
process (clock_c) begin
  if rising_edge(clock_c) then
    if i5 = "1" then
      n13 <= "0";
    elsif i4 = "1" then
      n13 <= n12;
    end if;
  end if;
end process;
process (clock_c) begin
  if rising_edge(clock_c) then
    if i5 = "1" then
      n14 <= "0";
    elsif i4 = "1" then
      n14 <= n13;
    end if;
  end if;
end process;
process (clock_c) begin
  if rising_edge(clock_c) then
    if i5 = "1" then
      n15 <= "0";
    elsif i4 = "1" then
      n15 <= n14;
    end if;
  end if;
end process;
process (clock_c) begin
  if rising_edge(clock_c) then
    if i5 = "1" then
      n16 <= "0";
    elsif i4 = "1" then
      n16 <= n15;
    end if;
  end if;
end process;
n17 <= not n16;
n18 <= s28_2 & s28_1;
n19 <= s28_3(31 downto 31) &
  s28_3(30 downto 30) &
  s28_3(29 downto 29) &
  s28_3(28 downto 28) &
  s28_3(27 downto 27) &
  s28_3(26 downto 26) &
  s28_3(25 downto 25) &
  s28_3(24 downto 24) &
  s28_3(23 downto 23) &
  s28_3(22 downto 22) &
  s28_3(21 downto 21) &
  s28_3(20 downto 20) &
  s28_3(19 downto 19) &
  s28_3(18 downto 18) &
  s28_3(17 downto 17) &
  s28_3(16 downto 16);
n20 <= s28_3(15 downto 15) &
  s28_3(14 downto 14) &
  s28_3(13 downto 13) &
  s28_3(12 downto 12) &
  s28_3(11 downto 11) &
  s28_3(10 downto 10) &
  s28_3(9 downto 9) &
  s28_3(8 downto 8) &
  s28_3(7 downto 7) &
  s28_3(6 downto 6) &
  s28_3(5 downto 5) &
  s28_3(4 downto 4) &
  s28_3(3 downto 3) &
  s28_3(2 downto 2) &
  s28_3(1 downto 1) &
  s28_3(0 downto 0);
n21 <= s29_1(31 downto 31) &
  s29_1(30 downto 30) &
  s29_1(29 downto 29) &
  s29_1(28 downto 28) &
  s29_1(27 downto 27) &
  s29_1(26 downto 26) &
  s29_1(25 downto 25) &
  s29_1(24 downto 24) &
  s29_1(23 downto 23) &
  s29_1(22 downto 22) &
  s29_1(21 downto 21) &
  s29_1(20 downto 20) &
  s29_1(19 downto 19) &
  s29_1(18 downto 18) &
  s29_1(17 downto 17) &
  s29_1(16 downto 16);
n22 <= s29_1(15 downto 15) &
  s29_1(14 downto 14) &
  s29_1(13 downto 13) &
  s29_1(12 downto 12) &
  s29_1(11 downto 11) &
  s29_1(10 downto 10) &
  s29_1(9 downto 9) &
  s29_1(8 downto 8) &
  s29_1(7 downto 7) &
  s29_1(6 downto 6) &
  s29_1(5 downto 5) &
  s29_1(4 downto 4) &
  s29_1(3 downto 3) &
  s29_1(2 downto 2) &
  s29_1(1 downto 1) &
  s29_1(0 downto 0);
n23 <= n20 when s25_1 = "1" else n19;
n24 <= n22 when s25_1 = "1" else n21;
s25 : cf_fft_2048_8_35 port map (clock_c, n18, i4, i5, s25_1);
s26 : cf_fft_2048_8_14 port map (clock_c, i2, i3, n1, i4, i5, s26_1, s26_2);
s27 : cf_fft_2048_8_26 port map (clock_c, i1, i4, i5, s27_1, s27_2);
s28 : cf_fft_2048_8_30 port map (clock_c, n2, n6, n11, n17, i4, i5, s28_1, s28_2, s28_3);
s29 : cf_fft_2048_8_31 port map (clock_c, n2, n6, n11, n16, i4, i5, s29_1);
o3 <= n24;
o2 <= n23;
o1 <= s28_1;
end architecture rtl;

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
entity cf_fft_2048_8_12 is
port (
clock_c : in std_logic;
i1 : in  unsigned(15 downto 0);
i2 : in  unsigned(15 downto 0);
i3 : in  unsigned(3 downto 0);
i4 : in  unsigned(0 downto 0);
i5 : in  unsigned(0 downto 0);
o1 : out unsigned(15 downto 0);
o2 : out unsigned(15 downto 0));
end entity cf_fft_2048_8_12;
architecture rtl of cf_fft_2048_8_12 is
signal n1 : unsigned(15 downto 0) := "0000000000000000";
signal n2 : unsigned(7 downto 0);
signal n3 : unsigned(7 downto 0);
signal n4 : unsigned(15 downto 0) := "0000000000000000";
signal n5 : unsigned(7 downto 0);
signal n6 : unsigned(7 downto 0);
signal n7 : unsigned(7 downto 0) := "00000000";
signal n8 : unsigned(7 downto 0) := "00000000";
signal n9 : unsigned(7 downto 0) := "00000000";
signal n10 : unsigned(7 downto 0) := "00000000";
signal n11 : unsigned(15 downto 0) := "0000000000000000";
signal n12 : unsigned(7 downto 0);
signal n13 : unsigned(7 downto 0);
signal n14 : unsigned(15 downto 0);
signal n15 : unsigned(7 downto 0);
signal n16 : unsigned(7 downto 0) := "00000000";
signal n17 : unsigned(15 downto 0);
signal n18 : unsigned(7 downto 0);
signal n19 : unsigned(7 downto 0) := "00000000";
signal n20 : unsigned(7 downto 0);
signal n21 : unsigned(7 downto 0) := "00000000";
signal n22 : unsigned(15 downto 0);
signal n23 : unsigned(7 downto 0);
signal n24 : unsigned(7 downto 0) := "00000000";
signal n25 : unsigned(15 downto 0);
signal n26 : unsigned(7 downto 0);
signal n27 : unsigned(7 downto 0) := "00000000";
signal n28 : unsigned(7 downto 0);
signal n29 : unsigned(7 downto 0) := "00000000";
signal n30 : unsigned(7 downto 0);
signal n31 : unsigned(7 downto 0);
signal n32 : unsigned(15 downto 0);
signal n33 : unsigned(15 downto 0) := "0000000000000000";
signal n34 : unsigned(7 downto 0);
signal n35 : unsigned(7 downto 0);
signal n36 : unsigned(15 downto 0);
signal n37 : unsigned(15 downto 0) := "0000000000000000";
begin
process (clock_c) begin
  if rising_edge(clock_c) then
    if i5 = "1" then
      n1 <= "0000000000000000";
    elsif i4 = "1" then
      n1 <= i1;
    end if;
  end if;
end process;
n2 <= n1(15 downto 15) &
  n1(14 downto 14) &
  n1(13 downto 13) &
  n1(12 downto 12) &
  n1(11 downto 11) &
  n1(10 downto 10) &
  n1(9 downto 9) &
  n1(8 downto 8);
n3 <= n1(7 downto 7) &
  n1(6 downto 6) &
  n1(5 downto 5) &
  n1(4 downto 4) &
  n1(3 downto 3) &
  n1(2 downto 2) &
  n1(1 downto 1) &
  n1(0 downto 0);
process (clock_c) begin
  if rising_edge(clock_c) then
    if i5 = "1" then
      n4 <= "0000000000000000";
    elsif i4 = "1" then
      n4 <= i2;
    end if;
  end if;
end process;
n5 <= n4(15 downto 15) &
  n4(14 downto 14) &
  n4(13 downto 13) &
  n4(12 downto 12) &
  n4(11 downto 11) &
  n4(10 downto 10) &
  n4(9 downto 9) &
  n4(8 downto 8);
n6 <= n4(7 downto 7) &
  n4(6 downto 6) &
  n4(5 downto 5) &
  n4(4 downto 4) &
  n4(3 downto 3) &
  n4(2 downto 2) &
  n4(1 downto 1) &
  n4(0 downto 0);
process (clock_c) begin
  if rising_edge(clock_c) then
    if i5 = "1" then
      n7 <= "00000000";
    elsif i4 = "1" then
      n7 <= n2;
    end if;
  end if;
end process;
process (clock_c) begin
  if rising_edge(clock_c) then
    if i5 = "1" then
      n8 <= "00000000";
    elsif i4 = "1" then
      n8 <= n7;
    end if;
  end if;
end process;
process (clock_c) begin
  if rising_edge(clock_c) then
    if i5 = "1" then
      n9 <= "00000000";
    elsif i4 = "1" then
      n9 <= n3;
    end if;
  end if;
end process;
process (clock_c) begin
  if rising_edge(clock_c) then
    if i5 = "1" then
      n10 <= "00000000";
    elsif i4 = "1" then
      n10 <= n9;
    end if;
  end if;
end process;
process (clock_c) begin
  if rising_edge(clock_c) then 
    if i4 = "1" then
      case i3 is
        when "0000" => n11 <= "0111111100000000";
        when "0001" => n11 <= "0111110111100111";
        when "0010" => n11 <= "0111011011001111";
        when "0011" => n11 <= "0110101010111000";
        when "0100" => n11 <= "0101101010100101";
        when "0101" => n11 <= "0100011110010101";
        when "0110" => n11 <= "0011000010001001";
        when "0111" => n11 <= "0001100010000010";
        when "1000" => n11 <= "0000000010000000";
        when "1001" => n11 <= "1110011110000010";
        when "1010" => n11 <= "1100111110001001";
        when "1011" => n11 <= "1011100010010101";
        when "1100" => n11 <= "1010010110100101";
        when "1101" => n11 <= "1001010110111000";
        when "1110" => n11 <= "1000100111001111";
        when "1111" => n11 <= "1000001011100111";
        when others => n11 <= "XXXXXXXXXXXXXXXX";
      end case;
    end if;
  end if;
end process;
n12 <= n11(15 downto 15) &
  n11(14 downto 14) &
  n11(13 downto 13) &
  n11(12 downto 12) &
  n11(11 downto 11) &
  n11(10 downto 10) &
  n11(9 downto 9) &
  n11(8 downto 8);
n13 <= n11(7 downto 7) &
  n11(6 downto 6) &
  n11(5 downto 5) &
  n11(4 downto 4) &
  n11(3 downto 3) &
  n11(2 downto 2) &
  n11(1 downto 1) &
  n11(0 downto 0);
n14 <= unsigned(signed(n5) * signed(n12));
n15 <= n14(14 downto 14) &
  n14(13 downto 13) &
  n14(12 downto 12) &
  n14(11 downto 11) &
  n14(10 downto 10) &
  n14(9 downto 9) &
  n14(8 downto 8) &
  n14(7 downto 7);
process (clock_c) begin
  if rising_edge(clock_c) then
    if i5 = "1" then
      n16 <= "00000000";
    elsif i4 = "1" then
      n16 <= n15;
    end if;
  end if;
end process;
n17 <= unsigned(signed(n6) * signed(n13));
n18 <= n17(14 downto 14) &
  n17(13 downto 13) &
  n17(12 downto 12) &
  n17(11 downto 11) &
  n17(10 downto 10) &
  n17(9 downto 9) &
  n17(8 downto 8) &
  n17(7 downto 7);
process (clock_c) begin
  if rising_edge(clock_c) then
    if i5 = "1" then
      n19 <= "00000000";
    elsif i4 = "1" then
      n19 <= n18;
    end if;
  end if;
end process;
n20 <= n16 - n19;
process (clock_c) begin
  if rising_edge(clock_c) then
    if i5 = "1" then
      n21 <= "00000000";
    elsif i4 = "1" then
      n21 <= n20;
    end if;
  end if;
end process;
n22 <= unsigned(signed(n5) * signed(n13));
n23 <= n22(14 downto 14) &
  n22(13 downto 13) &
  n22(12 downto 12) &
  n22(11 downto 11) &
  n22(10 downto 10) &
  n22(9 downto 9) &
  n22(8 downto 8) &
  n22(7 downto 7);
process (clock_c) begin
  if rising_edge(clock_c) then
    if i5 = "1" then
      n24 <= "00000000";
    elsif i4 = "1" then
      n24 <= n23;
    end if;
  end if;
end process;
n25 <= unsigned(signed(n6) * signed(n12));
n26 <= n25(14 downto 14) &
  n25(13 downto 13) &
  n25(12 downto 12) &
  n25(11 downto 11) &
  n25(10 downto 10) &
  n25(9 downto 9) &
  n25(8 downto 8) &
  n25(7 downto 7);
process (clock_c) begin
  if rising_edge(clock_c) then
    if i5 = "1" then
      n27 <= "00000000";
    elsif i4 = "1" then
      n27 <= n26;
    end if;
  end if;
end process;
n28 <= n24 + n27;
process (clock_c) begin
  if rising_edge(clock_c) then
    if i5 = "1" then
      n29 <= "00000000";
    elsif i4 = "1" then
      n29 <= n28;
    end if;
  end if;
end process;
n30 <= n8 + n21;
n31 <= n10 + n29;
n32 <= n30 & n31;
process (clock_c) begin
  if rising_edge(clock_c) then
    if i5 = "1" then
      n33 <= "0000000000000000";
    elsif i4 = "1" then
      n33 <= n32;
    end if;
  end if;
end process;
n34 <= n8 - n21;
n35 <= n10 - n29;
n36 <= n34 & n35;
process (clock_c) begin
  if rising_edge(clock_c) then
    if i5 = "1" then
      n37 <= "0000000000000000";
    elsif i4 = "1" then
      n37 <= n36;
    end if;
  end if;
end process;
o2 <= n37;
o1 <= n33;
end architecture rtl;

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
entity cf_fft_2048_8_11 is
port (
clock_c : in std_logic;
i1 : in  unsigned(0 downto 0);
i2 : in  unsigned(15 downto 0);
i3 : in  unsigned(15 downto 0);
i4 : in  unsigned(0 downto 0);
i5 : in  unsigned(0 downto 0);
o1 : out unsigned(0 downto 0);
o2 : out unsigned(15 downto 0);
o3 : out unsigned(15 downto 0));
end entity cf_fft_2048_8_11;
architecture rtl of cf_fft_2048_8_11 is
signal n1 : unsigned(3 downto 0);
signal n2 : unsigned(31 downto 0);
signal n3 : unsigned(0 downto 0) := "0";
signal n4 : unsigned(0 downto 0) := "0";
signal n5 : unsigned(0 downto 0) := "0";
signal n6 : unsigned(0 downto 0) := "0";
signal n7 : unsigned(8 downto 0);
signal n8 : unsigned(8 downto 0) := "000000000";
signal n9 : unsigned(8 downto 0) := "000000000";
signal n10 : unsigned(8 downto 0) := "000000000";
signal n11 : unsigned(8 downto 0) := "000000000";
signal n12 : unsigned(0 downto 0);
signal n13 : unsigned(0 downto 0) := "0";
signal n14 : unsigned(0 downto 0) := "0";
signal n15 : unsigned(0 downto 0) := "0";
signal n16 : unsigned(0 downto 0) := "0";
signal n17 : unsigned(0 downto 0);
signal n18 : unsigned(1 downto 0);
signal n19 : unsigned(15 downto 0);
signal n20 : unsigned(15 downto 0);
signal n21 : unsigned(15 downto 0);
signal n22 : unsigned(15 downto 0);
signal n23 : unsigned(15 downto 0);
signal n24 : unsigned(15 downto 0);
signal s25_1 : unsigned(0 downto 0);
signal s26_1 : unsigned(15 downto 0);
signal s26_2 : unsigned(15 downto 0);
signal s27_1 : unsigned(9 downto 0);
signal s27_2 : unsigned(0 downto 0);
signal s28_1 : unsigned(0 downto 0);
signal s28_2 : unsigned(0 downto 0);
signal s28_3 : unsigned(31 downto 0);
signal s29_1 : unsigned(31 downto 0);
component cf_fft_2048_8_35 is
port (
clock_c : in std_logic;
i1 : in  unsigned(1 downto 0);
i2 : in  unsigned(0 downto 0);
i3 : in  unsigned(0 downto 0);
o1 : out unsigned(0 downto 0));
end component cf_fft_2048_8_35;
component cf_fft_2048_8_12 is
port (
clock_c : in std_logic;
i1 : in  unsigned(15 downto 0);
i2 : in  unsigned(15 downto 0);
i3 : in  unsigned(3 downto 0);
i4 : in  unsigned(0 downto 0);
i5 : in  unsigned(0 downto 0);
o1 : out unsigned(15 downto 0);
o2 : out unsigned(15 downto 0));
end component cf_fft_2048_8_12;
component cf_fft_2048_8_26 is
port (
clock_c : in std_logic;
i1 : in  unsigned(0 downto 0);
i2 : in  unsigned(0 downto 0);
i3 : in  unsigned(0 downto 0);
o1 : out unsigned(9 downto 0);
o2 : out unsigned(0 downto 0));
end component cf_fft_2048_8_26;
component cf_fft_2048_8_30 is
port (
clock_c : in std_logic;
i1 : in  unsigned(31 downto 0);
i2 : in  unsigned(0 downto 0);
i3 : in  unsigned(8 downto 0);
i4 : in  unsigned(0 downto 0);
i5 : in  unsigned(0 downto 0);
i6 : in  unsigned(0 downto 0);
o1 : out unsigned(0 downto 0);
o2 : out unsigned(0 downto 0);
o3 : out unsigned(31 downto 0));
end component cf_fft_2048_8_30;
component cf_fft_2048_8_31 is
port (
clock_c : in std_logic;
i1 : in  unsigned(31 downto 0);
i2 : in  unsigned(0 downto 0);
i3 : in  unsigned(8 downto 0);
i4 : in  unsigned(0 downto 0);
i5 : in  unsigned(0 downto 0);
i6 : in  unsigned(0 downto 0);
o1 : out unsigned(31 downto 0));
end component cf_fft_2048_8_31;
begin
n1 <= s27_1(9 downto 9) &
  s27_1(8 downto 8) &
  s27_1(7 downto 7) &
  s27_1(6 downto 6);
n2 <= s26_1 & s26_2;
process (clock_c) begin
  if rising_edge(clock_c) then
    if i5 = "1" then
      n3 <= "0";
    elsif i4 = "1" then
      n3 <= s27_2;
    end if;
  end if;
end process;
process (clock_c) begin
  if rising_edge(clock_c) then
    if i5 = "1" then
      n4 <= "0";
    elsif i4 = "1" then
      n4 <= n3;
    end if;
  end if;
end process;
process (clock_c) begin
  if rising_edge(clock_c) then
    if i5 = "1" then
      n5 <= "0";
    elsif i4 = "1" then
      n5 <= n4;
    end if;
  end if;
end process;
process (clock_c) begin
  if rising_edge(clock_c) then
    if i5 = "1" then
      n6 <= "0";
    elsif i4 = "1" then
      n6 <= n5;
    end if;
  end if;
end process;
n7 <= s27_1(9 downto 9) &
  s27_1(8 downto 8) &
  s27_1(7 downto 7) &
  s27_1(6 downto 6) &
  s27_1(5 downto 5) &
  s27_1(4 downto 4) &
  s27_1(3 downto 3) &
  s27_1(2 downto 2) &
  s27_1(1 downto 1);
process (clock_c) begin
  if rising_edge(clock_c) then
    if i5 = "1" then
      n8 <= "000000000";
    elsif i4 = "1" then
      n8 <= n7;
    end if;
  end if;
end process;
process (clock_c) begin
  if rising_edge(clock_c) then
    if i5 = "1" then
      n9 <= "000000000";
    elsif i4 = "1" then
      n9 <= n8;
    end if;
  end if;
end process;
process (clock_c) begin
  if rising_edge(clock_c) then
    if i5 = "1" then
      n10 <= "000000000";
    elsif i4 = "1" then
      n10 <= n9;
    end if;
  end if;
end process;
process (clock_c) begin
  if rising_edge(clock_c) then
    if i5 = "1" then
      n11 <= "000000000";
    elsif i4 = "1" then
      n11 <= n10;
    end if;
  end if;
end process;
n12 <= s27_1(0 downto 0);
process (clock_c) begin
  if rising_edge(clock_c) then
    if i5 = "1" then
      n13 <= "0";
    elsif i4 = "1" then
      n13 <= n12;
    end if;
  end if;
end process;
process (clock_c) begin
  if rising_edge(clock_c) then
    if i5 = "1" then
      n14 <= "0";
    elsif i4 = "1" then
      n14 <= n13;
    end if;
  end if;
end process;
process (clock_c) begin
  if rising_edge(clock_c) then
    if i5 = "1" then
      n15 <= "0";
    elsif i4 = "1" then
      n15 <= n14;
    end if;
  end if;
end process;
process (clock_c) begin
  if rising_edge(clock_c) then
    if i5 = "1" then
      n16 <= "0";
    elsif i4 = "1" then
      n16 <= n15;
    end if;
  end if;
end process;
n17 <= not n16;
n18 <= s28_2 & s28_1;
n19 <= s28_3(31 downto 31) &
  s28_3(30 downto 30) &
  s28_3(29 downto 29) &
  s28_3(28 downto 28) &
  s28_3(27 downto 27) &
  s28_3(26 downto 26) &
  s28_3(25 downto 25) &
  s28_3(24 downto 24) &
  s28_3(23 downto 23) &
  s28_3(22 downto 22) &
  s28_3(21 downto 21) &
  s28_3(20 downto 20) &
  s28_3(19 downto 19) &
  s28_3(18 downto 18) &
  s28_3(17 downto 17) &
  s28_3(16 downto 16);
n20 <= s28_3(15 downto 15) &
  s28_3(14 downto 14) &
  s28_3(13 downto 13) &
  s28_3(12 downto 12) &
  s28_3(11 downto 11) &
  s28_3(10 downto 10) &
  s28_3(9 downto 9) &
  s28_3(8 downto 8) &
  s28_3(7 downto 7) &
  s28_3(6 downto 6) &
  s28_3(5 downto 5) &
  s28_3(4 downto 4) &
  s28_3(3 downto 3) &
  s28_3(2 downto 2) &
  s28_3(1 downto 1) &
  s28_3(0 downto 0);
n21 <= s29_1(31 downto 31) &
  s29_1(30 downto 30) &
  s29_1(29 downto 29) &
  s29_1(28 downto 28) &
  s29_1(27 downto 27) &
  s29_1(26 downto 26) &
  s29_1(25 downto 25) &
  s29_1(24 downto 24) &
  s29_1(23 downto 23) &
  s29_1(22 downto 22) &
  s29_1(21 downto 21) &
  s29_1(20 downto 20) &
  s29_1(19 downto 19) &
  s29_1(18 downto 18) &
  s29_1(17 downto 17) &
  s29_1(16 downto 16);
n22 <= s29_1(15 downto 15) &
  s29_1(14 downto 14) &
  s29_1(13 downto 13) &
  s29_1(12 downto 12) &
  s29_1(11 downto 11) &
  s29_1(10 downto 10) &
  s29_1(9 downto 9) &
  s29_1(8 downto 8) &
  s29_1(7 downto 7) &
  s29_1(6 downto 6) &
  s29_1(5 downto 5) &
  s29_1(4 downto 4) &
  s29_1(3 downto 3) &
  s29_1(2 downto 2) &
  s29_1(1 downto 1) &
  s29_1(0 downto 0);
n23 <= n20 when s25_1 = "1" else n19;
n24 <= n22 when s25_1 = "1" else n21;
s25 : cf_fft_2048_8_35 port map (clock_c, n18, i4, i5, s25_1);
s26 : cf_fft_2048_8_12 port map (clock_c, i2, i3, n1, i4, i5, s26_1, s26_2);
s27 : cf_fft_2048_8_26 port map (clock_c, i1, i4, i5, s27_1, s27_2);
s28 : cf_fft_2048_8_30 port map (clock_c, n2, n6, n11, n17, i4, i5, s28_1, s28_2, s28_3);
s29 : cf_fft_2048_8_31 port map (clock_c, n2, n6, n11, n16, i4, i5, s29_1);
o3 <= n24;
o2 <= n23;
o1 <= s28_1;
end architecture rtl;

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
entity cf_fft_2048_8_10 is
port (
clock_c : in std_logic;
i1 : in  unsigned(15 downto 0);
i2 : in  unsigned(15 downto 0);
i3 : in  unsigned(2 downto 0);
i4 : in  unsigned(0 downto 0);
i5 : in  unsigned(0 downto 0);
o1 : out unsigned(15 downto 0);
o2 : out unsigned(15 downto 0));
end entity cf_fft_2048_8_10;
architecture rtl of cf_fft_2048_8_10 is
signal n1 : unsigned(15 downto 0) := "0000000000000000";
signal n2 : unsigned(7 downto 0);
signal n3 : unsigned(7 downto 0);
signal n4 : unsigned(15 downto 0) := "0000000000000000";
signal n5 : unsigned(7 downto 0);
signal n6 : unsigned(7 downto 0);
signal n7 : unsigned(7 downto 0) := "00000000";
signal n8 : unsigned(7 downto 0) := "00000000";
signal n9 : unsigned(7 downto 0) := "00000000";
signal n10 : unsigned(7 downto 0) := "00000000";
signal n11 : unsigned(15 downto 0) := "0000000000000000";
signal n12 : unsigned(7 downto 0);
signal n13 : unsigned(7 downto 0);
signal n14 : unsigned(15 downto 0);
signal n15 : unsigned(7 downto 0);
signal n16 : unsigned(7 downto 0) := "00000000";
signal n17 : unsigned(15 downto 0);
signal n18 : unsigned(7 downto 0);
signal n19 : unsigned(7 downto 0) := "00000000";
signal n20 : unsigned(7 downto 0);
signal n21 : unsigned(7 downto 0) := "00000000";
signal n22 : unsigned(15 downto 0);
signal n23 : unsigned(7 downto 0);
signal n24 : unsigned(7 downto 0) := "00000000";
signal n25 : unsigned(15 downto 0);
signal n26 : unsigned(7 downto 0);
signal n27 : unsigned(7 downto 0) := "00000000";
signal n28 : unsigned(7 downto 0);
signal n29 : unsigned(7 downto 0) := "00000000";
signal n30 : unsigned(7 downto 0);
signal n31 : unsigned(7 downto 0);
signal n32 : unsigned(15 downto 0);
signal n33 : unsigned(15 downto 0) := "0000000000000000";
signal n34 : unsigned(7 downto 0);
signal n35 : unsigned(7 downto 0);
signal n36 : unsigned(15 downto 0);
signal n37 : unsigned(15 downto 0) := "0000000000000000";
begin
process (clock_c) begin
  if rising_edge(clock_c) then
    if i5 = "1" then
      n1 <= "0000000000000000";
    elsif i4 = "1" then
      n1 <= i1;
    end if;
  end if;
end process;
n2 <= n1(15 downto 15) &
  n1(14 downto 14) &
  n1(13 downto 13) &
  n1(12 downto 12) &
  n1(11 downto 11) &
  n1(10 downto 10) &
  n1(9 downto 9) &
  n1(8 downto 8);
n3 <= n1(7 downto 7) &
  n1(6 downto 6) &
  n1(5 downto 5) &
  n1(4 downto 4) &
  n1(3 downto 3) &
  n1(2 downto 2) &
  n1(1 downto 1) &
  n1(0 downto 0);
process (clock_c) begin
  if rising_edge(clock_c) then
    if i5 = "1" then
      n4 <= "0000000000000000";
    elsif i4 = "1" then
      n4 <= i2;
    end if;
  end if;
end process;
n5 <= n4(15 downto 15) &
  n4(14 downto 14) &
  n4(13 downto 13) &
  n4(12 downto 12) &
  n4(11 downto 11) &
  n4(10 downto 10) &
  n4(9 downto 9) &
  n4(8 downto 8);
n6 <= n4(7 downto 7) &
  n4(6 downto 6) &
  n4(5 downto 5) &
  n4(4 downto 4) &
  n4(3 downto 3) &
  n4(2 downto 2) &
  n4(1 downto 1) &
  n4(0 downto 0);
process (clock_c) begin
  if rising_edge(clock_c) then
    if i5 = "1" then
      n7 <= "00000000";
    elsif i4 = "1" then
      n7 <= n2;
    end if;
  end if;
end process;
process (clock_c) begin
  if rising_edge(clock_c) then
    if i5 = "1" then
      n8 <= "00000000";
    elsif i4 = "1" then
      n8 <= n7;
    end if;
  end if;
end process;
process (clock_c) begin
  if rising_edge(clock_c) then
    if i5 = "1" then
      n9 <= "00000000";
    elsif i4 = "1" then
      n9 <= n3;
    end if;
  end if;
end process;
process (clock_c) begin
  if rising_edge(clock_c) then
    if i5 = "1" then
      n10 <= "00000000";
    elsif i4 = "1" then
      n10 <= n9;
    end if;
  end if;
end process;
process (clock_c) begin
  if rising_edge(clock_c) then 
    if i4 = "1" then
      case i3 is
        when "000" => n11 <= "0111111100000000";
        when "001" => n11 <= "0111011011001111";
        when "010" => n11 <= "0101101010100101";
        when "011" => n11 <= "0011000010001001";
        when "100" => n11 <= "0000000010000000";
        when "101" => n11 <= "1100111110001001";
        when "110" => n11 <= "1010010110100101";
        when "111" => n11 <= "1000100111001111";
        when others => n11 <= "XXXXXXXXXXXXXXXX";
      end case;
    end if;
  end if;
end process;
n12 <= n11(15 downto 15) &
  n11(14 downto 14) &
  n11(13 downto 13) &
  n11(12 downto 12) &
  n11(11 downto 11) &
  n11(10 downto 10) &
  n11(9 downto 9) &
  n11(8 downto 8);
n13 <= n11(7 downto 7) &
  n11(6 downto 6) &
  n11(5 downto 5) &
  n11(4 downto 4) &
  n11(3 downto 3) &
  n11(2 downto 2) &
  n11(1 downto 1) &
  n11(0 downto 0);
n14 <= unsigned(signed(n5) * signed(n12));
n15 <= n14(14 downto 14) &
  n14(13 downto 13) &
  n14(12 downto 12) &
  n14(11 downto 11) &
  n14(10 downto 10) &
  n14(9 downto 9) &
  n14(8 downto 8) &
  n14(7 downto 7);
process (clock_c) begin
  if rising_edge(clock_c) then
    if i5 = "1" then
      n16 <= "00000000";
    elsif i4 = "1" then
      n16 <= n15;
    end if;
  end if;
end process;
n17 <= unsigned(signed(n6) * signed(n13));
n18 <= n17(14 downto 14) &
  n17(13 downto 13) &
  n17(12 downto 12) &
  n17(11 downto 11) &
  n17(10 downto 10) &
  n17(9 downto 9) &
  n17(8 downto 8) &
  n17(7 downto 7);
process (clock_c) begin
  if rising_edge(clock_c) then
    if i5 = "1" then
      n19 <= "00000000";
    elsif i4 = "1" then
      n19 <= n18;
    end if;
  end if;
end process;
n20 <= n16 - n19;
process (clock_c) begin
  if rising_edge(clock_c) then
    if i5 = "1" then
      n21 <= "00000000";
    elsif i4 = "1" then
      n21 <= n20;
    end if;
  end if;
end process;
n22 <= unsigned(signed(n5) * signed(n13));
n23 <= n22(14 downto 14) &
  n22(13 downto 13) &
  n22(12 downto 12) &
  n22(11 downto 11) &
  n22(10 downto 10) &
  n22(9 downto 9) &
  n22(8 downto 8) &
  n22(7 downto 7);
process (clock_c) begin
  if rising_edge(clock_c) then
    if i5 = "1" then
      n24 <= "00000000";
    elsif i4 = "1" then
      n24 <= n23;
    end if;
  end if;
end process;
n25 <= unsigned(signed(n6) * signed(n12));
n26 <= n25(14 downto 14) &
  n25(13 downto 13) &
  n25(12 downto 12) &
  n25(11 downto 11) &
  n25(10 downto 10) &
  n25(9 downto 9) &
  n25(8 downto 8) &
  n25(7 downto 7);
process (clock_c) begin
  if rising_edge(clock_c) then
    if i5 = "1" then
      n27 <= "00000000";
    elsif i4 = "1" then
      n27 <= n26;
    end if;
  end if;
end process;
n28 <= n24 + n27;
process (clock_c) begin
  if rising_edge(clock_c) then
    if i5 = "1" then
      n29 <= "00000000";
    elsif i4 = "1" then
      n29 <= n28;
    end if;
  end if;
end process;
n30 <= n8 + n21;
n31 <= n10 + n29;
n32 <= n30 & n31;
process (clock_c) begin
  if rising_edge(clock_c) then
    if i5 = "1" then
      n33 <= "0000000000000000";
    elsif i4 = "1" then
      n33 <= n32;
    end if;
  end if;
end process;
n34 <= n8 - n21;
n35 <= n10 - n29;
n36 <= n34 & n35;
process (clock_c) begin
  if rising_edge(clock_c) then
    if i5 = "1" then
      n37 <= "0000000000000000";
    elsif i4 = "1" then
      n37 <= n36;
    end if;
  end if;
end process;
o2 <= n37;
o1 <= n33;
end architecture rtl;

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
entity cf_fft_2048_8_9 is
port (
clock_c : in std_logic;
i1 : in  unsigned(0 downto 0);
i2 : in  unsigned(15 downto 0);
i3 : in  unsigned(15 downto 0);
i4 : in  unsigned(0 downto 0);
i5 : in  unsigned(0 downto 0);
o1 : out unsigned(0 downto 0);
o2 : out unsigned(15 downto 0);
o3 : out unsigned(15 downto 0));
end entity cf_fft_2048_8_9;
architecture rtl of cf_fft_2048_8_9 is
signal n1 : unsigned(2 downto 0);
signal n2 : unsigned(31 downto 0);
signal n3 : unsigned(0 downto 0) := "0";
signal n4 : unsigned(0 downto 0) := "0";
signal n5 : unsigned(0 downto 0) := "0";
signal n6 : unsigned(0 downto 0) := "0";
signal n7 : unsigned(8 downto 0);
signal n8 : unsigned(8 downto 0) := "000000000";
signal n9 : unsigned(8 downto 0) := "000000000";
signal n10 : unsigned(8 downto 0) := "000000000";
signal n11 : unsigned(8 downto 0) := "000000000";
signal n12 : unsigned(0 downto 0);
signal n13 : unsigned(0 downto 0) := "0";
signal n14 : unsigned(0 downto 0) := "0";
signal n15 : unsigned(0 downto 0) := "0";
signal n16 : unsigned(0 downto 0) := "0";
signal n17 : unsigned(0 downto 0);
signal n18 : unsigned(1 downto 0);
signal n19 : unsigned(15 downto 0);
signal n20 : unsigned(15 downto 0);
signal n21 : unsigned(15 downto 0);
signal n22 : unsigned(15 downto 0);
signal n23 : unsigned(15 downto 0);
signal n24 : unsigned(15 downto 0);
signal s25_1 : unsigned(15 downto 0);
signal s25_2 : unsigned(15 downto 0);
signal s26_1 : unsigned(0 downto 0);
signal s27_1 : unsigned(0 downto 0);
signal s27_2 : unsigned(0 downto 0);
signal s27_3 : unsigned(31 downto 0);
signal s28_1 : unsigned(31 downto 0);
signal s29_1 : unsigned(9 downto 0);
signal s29_2 : unsigned(0 downto 0);
component cf_fft_2048_8_10 is
port (
clock_c : in std_logic;
i1 : in  unsigned(15 downto 0);
i2 : in  unsigned(15 downto 0);
i3 : in  unsigned(2 downto 0);
i4 : in  unsigned(0 downto 0);
i5 : in  unsigned(0 downto 0);
o1 : out unsigned(15 downto 0);
o2 : out unsigned(15 downto 0));
end component cf_fft_2048_8_10;
component cf_fft_2048_8_35 is
port (
clock_c : in std_logic;
i1 : in  unsigned(1 downto 0);
i2 : in  unsigned(0 downto 0);
i3 : in  unsigned(0 downto 0);
o1 : out unsigned(0 downto 0));
end component cf_fft_2048_8_35;
component cf_fft_2048_8_30 is
port (
clock_c : in std_logic;
i1 : in  unsigned(31 downto 0);
i2 : in  unsigned(0 downto 0);
i3 : in  unsigned(8 downto 0);
i4 : in  unsigned(0 downto 0);
i5 : in  unsigned(0 downto 0);
i6 : in  unsigned(0 downto 0);
o1 : out unsigned(0 downto 0);
o2 : out unsigned(0 downto 0);
o3 : out unsigned(31 downto 0));
end component cf_fft_2048_8_30;
component cf_fft_2048_8_31 is
port (
clock_c : in std_logic;
i1 : in  unsigned(31 downto 0);
i2 : in  unsigned(0 downto 0);
i3 : in  unsigned(8 downto 0);
i4 : in  unsigned(0 downto 0);
i5 : in  unsigned(0 downto 0);
i6 : in  unsigned(0 downto 0);
o1 : out unsigned(31 downto 0));
end component cf_fft_2048_8_31;
component cf_fft_2048_8_26 is
port (
clock_c : in std_logic;
i1 : in  unsigned(0 downto 0);
i2 : in  unsigned(0 downto 0);
i3 : in  unsigned(0 downto 0);
o1 : out unsigned(9 downto 0);
o2 : out unsigned(0 downto 0));
end component cf_fft_2048_8_26;
begin
n1 <= s29_1(9 downto 9) &
  s29_1(8 downto 8) &
  s29_1(7 downto 7);
n2 <= s25_1 & s25_2;
process (clock_c) begin
  if rising_edge(clock_c) then
    if i5 = "1" then
      n3 <= "0";
    elsif i4 = "1" then
      n3 <= s29_2;
    end if;
  end if;
end process;
process (clock_c) begin
  if rising_edge(clock_c) then
    if i5 = "1" then
      n4 <= "0";
    elsif i4 = "1" then
      n4 <= n3;
    end if;
  end if;
end process;
process (clock_c) begin
  if rising_edge(clock_c) then
    if i5 = "1" then
      n5 <= "0";
    elsif i4 = "1" then
      n5 <= n4;
    end if;
  end if;
end process;
process (clock_c) begin
  if rising_edge(clock_c) then
    if i5 = "1" then
      n6 <= "0";
    elsif i4 = "1" then
      n6 <= n5;
    end if;
  end if;
end process;
n7 <= s29_1(9 downto 9) &
  s29_1(8 downto 8) &
  s29_1(7 downto 7) &
  s29_1(6 downto 6) &
  s29_1(5 downto 5) &
  s29_1(4 downto 4) &
  s29_1(3 downto 3) &
  s29_1(2 downto 2) &
  s29_1(1 downto 1);
process (clock_c) begin
  if rising_edge(clock_c) then
    if i5 = "1" then
      n8 <= "000000000";
    elsif i4 = "1" then
      n8 <= n7;
    end if;
  end if;
end process;
process (clock_c) begin
  if rising_edge(clock_c) then
    if i5 = "1" then
      n9 <= "000000000";
    elsif i4 = "1" then
      n9 <= n8;
    end if;
  end if;
end process;
process (clock_c) begin
  if rising_edge(clock_c) then
    if i5 = "1" then
      n10 <= "000000000";
    elsif i4 = "1" then
      n10 <= n9;
    end if;
  end if;
end process;
process (clock_c) begin
  if rising_edge(clock_c) then
    if i5 = "1" then
      n11 <= "000000000";
    elsif i4 = "1" then
      n11 <= n10;
    end if;
  end if;
end process;
n12 <= s29_1(0 downto 0);
process (clock_c) begin
  if rising_edge(clock_c) then
    if i5 = "1" then
      n13 <= "0";
    elsif i4 = "1" then
      n13 <= n12;
    end if;
  end if;
end process;
process (clock_c) begin
  if rising_edge(clock_c) then
    if i5 = "1" then
      n14 <= "0";
    elsif i4 = "1" then
      n14 <= n13;
    end if;
  end if;
end process;
process (clock_c) begin
  if rising_edge(clock_c) then
    if i5 = "1" then
      n15 <= "0";
    elsif i4 = "1" then
      n15 <= n14;
    end if;
  end if;
end process;
process (clock_c) begin
  if rising_edge(clock_c) then
    if i5 = "1" then
      n16 <= "0";
    elsif i4 = "1" then
      n16 <= n15;
    end if;
  end if;
end process;
n17 <= not n16;
n18 <= s27_2 & s27_1;
n19 <= s27_3(31 downto 31) &
  s27_3(30 downto 30) &
  s27_3(29 downto 29) &
  s27_3(28 downto 28) &
  s27_3(27 downto 27) &
  s27_3(26 downto 26) &
  s27_3(25 downto 25) &
  s27_3(24 downto 24) &
  s27_3(23 downto 23) &
  s27_3(22 downto 22) &
  s27_3(21 downto 21) &
  s27_3(20 downto 20) &
  s27_3(19 downto 19) &
  s27_3(18 downto 18) &
  s27_3(17 downto 17) &
  s27_3(16 downto 16);
n20 <= s27_3(15 downto 15) &
  s27_3(14 downto 14) &
  s27_3(13 downto 13) &
  s27_3(12 downto 12) &
  s27_3(11 downto 11) &
  s27_3(10 downto 10) &
  s27_3(9 downto 9) &
  s27_3(8 downto 8) &
  s27_3(7 downto 7) &
  s27_3(6 downto 6) &
  s27_3(5 downto 5) &
  s27_3(4 downto 4) &
  s27_3(3 downto 3) &
  s27_3(2 downto 2) &
  s27_3(1 downto 1) &
  s27_3(0 downto 0);
n21 <= s28_1(31 downto 31) &
  s28_1(30 downto 30) &
  s28_1(29 downto 29) &
  s28_1(28 downto 28) &
  s28_1(27 downto 27) &
  s28_1(26 downto 26) &
  s28_1(25 downto 25) &
  s28_1(24 downto 24) &
  s28_1(23 downto 23) &
  s28_1(22 downto 22) &
  s28_1(21 downto 21) &
  s28_1(20 downto 20) &
  s28_1(19 downto 19) &
  s28_1(18 downto 18) &
  s28_1(17 downto 17) &
  s28_1(16 downto 16);
n22 <= s28_1(15 downto 15) &
  s28_1(14 downto 14) &
  s28_1(13 downto 13) &
  s28_1(12 downto 12) &
  s28_1(11 downto 11) &
  s28_1(10 downto 10) &
  s28_1(9 downto 9) &
  s28_1(8 downto 8) &
  s28_1(7 downto 7) &
  s28_1(6 downto 6) &
  s28_1(5 downto 5) &
  s28_1(4 downto 4) &
  s28_1(3 downto 3) &
  s28_1(2 downto 2) &
  s28_1(1 downto 1) &
  s28_1(0 downto 0);
n23 <= n20 when s26_1 = "1" else n19;
n24 <= n22 when s26_1 = "1" else n21;
s25 : cf_fft_2048_8_10 port map (clock_c, i2, i3, n1, i4, i5, s25_1, s25_2);
s26 : cf_fft_2048_8_35 port map (clock_c, n18, i4, i5, s26_1);
s27 : cf_fft_2048_8_30 port map (clock_c, n2, n6, n11, n17, i4, i5, s27_1, s27_2, s27_3);
s28 : cf_fft_2048_8_31 port map (clock_c, n2, n6, n11, n16, i4, i5, s28_1);
s29 : cf_fft_2048_8_26 port map (clock_c, i1, i4, i5, s29_1, s29_2);
o3 <= n24;
o2 <= n23;
o1 <= s27_1;
end architecture rtl;

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
entity cf_fft_2048_8_8 is
port (
clock_c : in std_logic;
i1 : in  unsigned(0 downto 0);
i2 : in  unsigned(15 downto 0);
i3 : in  unsigned(15 downto 0);
i4 : in  unsigned(0 downto 0);
i5 : in  unsigned(0 downto 0);
o1 : out unsigned(0 downto 0);
o2 : out unsigned(15 downto 0);
o3 : out unsigned(15 downto 0));
end entity cf_fft_2048_8_8;
architecture rtl of cf_fft_2048_8_8 is
signal s1_1 : unsigned(0 downto 0);
signal s1_2 : unsigned(15 downto 0);
signal s1_3 : unsigned(15 downto 0);
signal s2_1 : unsigned(0 downto 0);
signal s2_2 : unsigned(15 downto 0);
signal s2_3 : unsigned(15 downto 0);
signal s3_1 : unsigned(0 downto 0);
signal s3_2 : unsigned(15 downto 0);
signal s3_3 : unsigned(15 downto 0);
signal s4_1 : unsigned(0 downto 0);
signal s4_2 : unsigned(15 downto 0);
signal s4_3 : unsigned(15 downto 0);
signal s5_1 : unsigned(0 downto 0);
signal s5_2 : unsigned(15 downto 0);
signal s5_3 : unsigned(15 downto 0);
signal s6_1 : unsigned(0 downto 0);
signal s6_2 : unsigned(15 downto 0);
signal s6_3 : unsigned(15 downto 0);
signal s7_1 : unsigned(0 downto 0);
signal s7_2 : unsigned(15 downto 0);
signal s7_3 : unsigned(15 downto 0);
signal s8_1 : unsigned(0 downto 0);
signal s8_2 : unsigned(15 downto 0);
signal s8_3 : unsigned(15 downto 0);
component cf_fft_2048_8_23 is
port (
clock_c : in std_logic;
i1 : in  unsigned(0 downto 0);
i2 : in  unsigned(15 downto 0);
i3 : in  unsigned(15 downto 0);
i4 : in  unsigned(0 downto 0);
i5 : in  unsigned(0 downto 0);
o1 : out unsigned(0 downto 0);
o2 : out unsigned(15 downto 0);
o3 : out unsigned(15 downto 0));
end component cf_fft_2048_8_23;
component cf_fft_2048_8_21 is
port (
clock_c : in std_logic;
i1 : in  unsigned(0 downto 0);
i2 : in  unsigned(15 downto 0);
i3 : in  unsigned(15 downto 0);
i4 : in  unsigned(0 downto 0);
i5 : in  unsigned(0 downto 0);
o1 : out unsigned(0 downto 0);
o2 : out unsigned(15 downto 0);
o3 : out unsigned(15 downto 0));
end component cf_fft_2048_8_21;
component cf_fft_2048_8_19 is
port (
clock_c : in std_logic;
i1 : in  unsigned(0 downto 0);
i2 : in  unsigned(15 downto 0);
i3 : in  unsigned(15 downto 0);
i4 : in  unsigned(0 downto 0);
i5 : in  unsigned(0 downto 0);
o1 : out unsigned(0 downto 0);
o2 : out unsigned(15 downto 0);
o3 : out unsigned(15 downto 0));
end component cf_fft_2048_8_19;
component cf_fft_2048_8_17 is
port (
clock_c : in std_logic;
i1 : in  unsigned(0 downto 0);
i2 : in  unsigned(15 downto 0);
i3 : in  unsigned(15 downto 0);
i4 : in  unsigned(0 downto 0);
i5 : in  unsigned(0 downto 0);
o1 : out unsigned(0 downto 0);
o2 : out unsigned(15 downto 0);
o3 : out unsigned(15 downto 0));
end component cf_fft_2048_8_17;
component cf_fft_2048_8_15 is
port (
clock_c : in std_logic;
i1 : in  unsigned(0 downto 0);
i2 : in  unsigned(15 downto 0);
i3 : in  unsigned(15 downto 0);
i4 : in  unsigned(0 downto 0);
i5 : in  unsigned(0 downto 0);
o1 : out unsigned(0 downto 0);
o2 : out unsigned(15 downto 0);
o3 : out unsigned(15 downto 0));
end component cf_fft_2048_8_15;
component cf_fft_2048_8_13 is
port (
clock_c : in std_logic;
i1 : in  unsigned(0 downto 0);
i2 : in  unsigned(15 downto 0);
i3 : in  unsigned(15 downto 0);
i4 : in  unsigned(0 downto 0);
i5 : in  unsigned(0 downto 0);
o1 : out unsigned(0 downto 0);
o2 : out unsigned(15 downto 0);
o3 : out unsigned(15 downto 0));
end component cf_fft_2048_8_13;
component cf_fft_2048_8_11 is
port (
clock_c : in std_logic;
i1 : in  unsigned(0 downto 0);
i2 : in  unsigned(15 downto 0);
i3 : in  unsigned(15 downto 0);
i4 : in  unsigned(0 downto 0);
i5 : in  unsigned(0 downto 0);
o1 : out unsigned(0 downto 0);
o2 : out unsigned(15 downto 0);
o3 : out unsigned(15 downto 0));
end component cf_fft_2048_8_11;
component cf_fft_2048_8_9 is
port (
clock_c : in std_logic;
i1 : in  unsigned(0 downto 0);
i2 : in  unsigned(15 downto 0);
i3 : in  unsigned(15 downto 0);
i4 : in  unsigned(0 downto 0);
i5 : in  unsigned(0 downto 0);
o1 : out unsigned(0 downto 0);
o2 : out unsigned(15 downto 0);
o3 : out unsigned(15 downto 0));
end component cf_fft_2048_8_9;
begin
s1 : cf_fft_2048_8_23 port map (clock_c, s2_1, s2_2, s2_3, i4, i5, s1_1, s1_2, s1_3);
s2 : cf_fft_2048_8_21 port map (clock_c, s3_1, s3_2, s3_3, i4, i5, s2_1, s2_2, s2_3);
s3 : cf_fft_2048_8_19 port map (clock_c, s4_1, s4_2, s4_3, i4, i5, s3_1, s3_2, s3_3);
s4 : cf_fft_2048_8_17 port map (clock_c, s5_1, s5_2, s5_3, i4, i5, s4_1, s4_2, s4_3);
s5 : cf_fft_2048_8_15 port map (clock_c, s6_1, s6_2, s6_3, i4, i5, s5_1, s5_2, s5_3);
s6 : cf_fft_2048_8_13 port map (clock_c, s7_1, s7_2, s7_3, i4, i5, s6_1, s6_2, s6_3);
s7 : cf_fft_2048_8_11 port map (clock_c, s8_1, s8_2, s8_3, i4, i5, s7_1, s7_2, s7_3);
s8 : cf_fft_2048_8_9 port map (clock_c, i1, i2, i3, i4, i5, s8_1, s8_2, s8_3);
o3 <= s1_3;
o2 <= s1_2;
o1 <= s1_1;
end architecture rtl;

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
entity cf_fft_2048_8_7 is
port (
clock_c : in std_logic;
i1 : in  unsigned(15 downto 0);
i2 : in  unsigned(15 downto 0);
i3 : in  unsigned(0 downto 0);
i4 : in  unsigned(0 downto 0);
i5 : in  unsigned(0 downto 0);
o1 : out unsigned(15 downto 0);
o2 : out unsigned(15 downto 0));
end entity cf_fft_2048_8_7;
architecture rtl of cf_fft_2048_8_7 is
signal n1 : unsigned(15 downto 0) := "0000000000000000";
signal n2 : unsigned(7 downto 0);
signal n3 : unsigned(7 downto 0);
signal n4 : unsigned(15 downto 0) := "0000000000000000";
signal n5 : unsigned(7 downto 0);
signal n6 : unsigned(7 downto 0);
signal n7 : unsigned(7 downto 0) := "00000000";
signal n8 : unsigned(7 downto 0) := "00000000";
signal n9 : unsigned(7 downto 0) := "00000000";
signal n10 : unsigned(7 downto 0) := "00000000";
signal n11 : unsigned(15 downto 0) := "0000000000000000";
signal n12 : unsigned(7 downto 0);
signal n13 : unsigned(7 downto 0);
signal n14 : unsigned(15 downto 0);
signal n15 : unsigned(7 downto 0);
signal n16 : unsigned(7 downto 0) := "00000000";
signal n17 : unsigned(15 downto 0);
signal n18 : unsigned(7 downto 0);
signal n19 : unsigned(7 downto 0) := "00000000";
signal n20 : unsigned(7 downto 0);
signal n21 : unsigned(7 downto 0) := "00000000";
signal n22 : unsigned(15 downto 0);
signal n23 : unsigned(7 downto 0);
signal n24 : unsigned(7 downto 0) := "00000000";
signal n25 : unsigned(15 downto 0);
signal n26 : unsigned(7 downto 0);
signal n27 : unsigned(7 downto 0) := "00000000";
signal n28 : unsigned(7 downto 0);
signal n29 : unsigned(7 downto 0) := "00000000";
signal n30 : unsigned(7 downto 0);
signal n31 : unsigned(7 downto 0);
signal n32 : unsigned(15 downto 0);
signal n33 : unsigned(15 downto 0) := "0000000000000000";
signal n34 : unsigned(7 downto 0);
signal n35 : unsigned(7 downto 0);
signal n36 : unsigned(15 downto 0);
signal n37 : unsigned(15 downto 0) := "0000000000000000";
begin
process (clock_c) begin
  if rising_edge(clock_c) then
    if i5 = "1" then
      n1 <= "0000000000000000";
    elsif i4 = "1" then
      n1 <= i1;
    end if;
  end if;
end process;
n2 <= n1(15 downto 15) &
  n1(14 downto 14) &
  n1(13 downto 13) &
  n1(12 downto 12) &
  n1(11 downto 11) &
  n1(10 downto 10) &
  n1(9 downto 9) &
  n1(8 downto 8);
n3 <= n1(7 downto 7) &
  n1(6 downto 6) &
  n1(5 downto 5) &
  n1(4 downto 4) &
  n1(3 downto 3) &
  n1(2 downto 2) &
  n1(1 downto 1) &
  n1(0 downto 0);
process (clock_c) begin
  if rising_edge(clock_c) then
    if i5 = "1" then
      n4 <= "0000000000000000";
    elsif i4 = "1" then
      n4 <= i2;
    end if;
  end if;
end process;
n5 <= n4(15 downto 15) &
  n4(14 downto 14) &
  n4(13 downto 13) &
  n4(12 downto 12) &
  n4(11 downto 11) &
  n4(10 downto 10) &
  n4(9 downto 9) &
  n4(8 downto 8);
n6 <= n4(7 downto 7) &
  n4(6 downto 6) &
  n4(5 downto 5) &
  n4(4 downto 4) &
  n4(3 downto 3) &
  n4(2 downto 2) &
  n4(1 downto 1) &
  n4(0 downto 0);
process (clock_c) begin
  if rising_edge(clock_c) then
    if i5 = "1" then
      n7 <= "00000000";
    elsif i4 = "1" then
      n7 <= n2;
    end if;
  end if;
end process;
process (clock_c) begin
  if rising_edge(clock_c) then
    if i5 = "1" then
      n8 <= "00000000";
    elsif i4 = "1" then
      n8 <= n7;
    end if;
  end if;
end process;
process (clock_c) begin
  if rising_edge(clock_c) then
    if i5 = "1" then
      n9 <= "00000000";
    elsif i4 = "1" then
      n9 <= n3;
    end if;
  end if;
end process;
process (clock_c) begin
  if rising_edge(clock_c) then
    if i5 = "1" then
      n10 <= "00000000";
    elsif i4 = "1" then
      n10 <= n9;
    end if;
  end if;
end process;
process (clock_c) begin
  if rising_edge(clock_c) then 
    if i4 = "1" then
      case i3 is
        when "0" => n11 <= "0111111100000000";
        when "1" => n11 <= "0000000010000000";
        when others => n11 <= "XXXXXXXXXXXXXXXX";
      end case;
    end if;
  end if;
end process;
n12 <= n11(15 downto 15) &
  n11(14 downto 14) &
  n11(13 downto 13) &
  n11(12 downto 12) &
  n11(11 downto 11) &
  n11(10 downto 10) &
  n11(9 downto 9) &
  n11(8 downto 8);
n13 <= n11(7 downto 7) &
  n11(6 downto 6) &
  n11(5 downto 5) &
  n11(4 downto 4) &
  n11(3 downto 3) &
  n11(2 downto 2) &
  n11(1 downto 1) &
  n11(0 downto 0);
n14 <= unsigned(signed(n5) * signed(n12));
n15 <= n14(14 downto 14) &
  n14(13 downto 13) &
  n14(12 downto 12) &
  n14(11 downto 11) &
  n14(10 downto 10) &
  n14(9 downto 9) &
  n14(8 downto 8) &
  n14(7 downto 7);
process (clock_c) begin
  if rising_edge(clock_c) then
    if i5 = "1" then
      n16 <= "00000000";
    elsif i4 = "1" then
      n16 <= n15;
    end if;
  end if;
end process;
n17 <= unsigned(signed(n6) * signed(n13));
n18 <= n17(14 downto 14) &
  n17(13 downto 13) &
  n17(12 downto 12) &
  n17(11 downto 11) &
  n17(10 downto 10) &
  n17(9 downto 9) &
  n17(8 downto 8) &
  n17(7 downto 7);
process (clock_c) begin
  if rising_edge(clock_c) then
    if i5 = "1" then
      n19 <= "00000000";
    elsif i4 = "1" then
      n19 <= n18;
    end if;
  end if;
end process;
n20 <= n16 - n19;
process (clock_c) begin
  if rising_edge(clock_c) then
    if i5 = "1" then
      n21 <= "00000000";
    elsif i4 = "1" then
      n21 <= n20;
    end if;
  end if;
end process;
n22 <= unsigned(signed(n5) * signed(n13));
n23 <= n22(14 downto 14) &
  n22(13 downto 13) &
  n22(12 downto 12) &
  n22(11 downto 11) &
  n22(10 downto 10) &
  n22(9 downto 9) &
  n22(8 downto 8) &
  n22(7 downto 7);
process (clock_c) begin
  if rising_edge(clock_c) then
    if i5 = "1" then
      n24 <= "00000000";
    elsif i4 = "1" then
      n24 <= n23;
    end if;
  end if;
end process;
n25 <= unsigned(signed(n6) * signed(n12));
n26 <= n25(14 downto 14) &
  n25(13 downto 13) &
  n25(12 downto 12) &
  n25(11 downto 11) &
  n25(10 downto 10) &
  n25(9 downto 9) &
  n25(8 downto 8) &
  n25(7 downto 7);
process (clock_c) begin
  if rising_edge(clock_c) then
    if i5 = "1" then
      n27 <= "00000000";
    elsif i4 = "1" then
      n27 <= n26;
    end if;
  end if;
end process;
n28 <= n24 + n27;
process (clock_c) begin
  if rising_edge(clock_c) then
    if i5 = "1" then
      n29 <= "00000000";
    elsif i4 = "1" then
      n29 <= n28;
    end if;
  end if;
end process;
n30 <= n8 + n21;
n31 <= n10 + n29;
n32 <= n30 & n31;
process (clock_c) begin
  if rising_edge(clock_c) then
    if i5 = "1" then
      n33 <= "0000000000000000";
    elsif i4 = "1" then
      n33 <= n32;
    end if;
  end if;
end process;
n34 <= n8 - n21;
n35 <= n10 - n29;
n36 <= n34 & n35;
process (clock_c) begin
  if rising_edge(clock_c) then
    if i5 = "1" then
      n37 <= "0000000000000000";
    elsif i4 = "1" then
      n37 <= n36;
    end if;
  end if;
end process;
o2 <= n37;
o1 <= n33;
end architecture rtl;

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
entity cf_fft_2048_8_6 is
port (
clock_c : in std_logic;
i1 : in  unsigned(0 downto 0);
i2 : in  unsigned(15 downto 0);
i3 : in  unsigned(15 downto 0);
i4 : in  unsigned(0 downto 0);
i5 : in  unsigned(0 downto 0);
o1 : out unsigned(0 downto 0);
o2 : out unsigned(15 downto 0);
o3 : out unsigned(15 downto 0));
end entity cf_fft_2048_8_6;
architecture rtl of cf_fft_2048_8_6 is
signal n1 : unsigned(0 downto 0);
signal n2 : unsigned(31 downto 0);
signal n3 : unsigned(0 downto 0) := "0";
signal n4 : unsigned(0 downto 0) := "0";
signal n5 : unsigned(0 downto 0) := "0";
signal n6 : unsigned(0 downto 0) := "0";
signal n7 : unsigned(8 downto 0);
signal n8 : unsigned(8 downto 0) := "000000000";
signal n9 : unsigned(8 downto 0) := "000000000";
signal n10 : unsigned(8 downto 0) := "000000000";
signal n11 : unsigned(8 downto 0) := "000000000";
signal n12 : unsigned(0 downto 0);
signal n13 : unsigned(0 downto 0) := "0";
signal n14 : unsigned(0 downto 0) := "0";
signal n15 : unsigned(0 downto 0) := "0";
signal n16 : unsigned(0 downto 0) := "0";
signal n17 : unsigned(0 downto 0);
signal n18 : unsigned(1 downto 0);
signal n19 : unsigned(15 downto 0);
signal n20 : unsigned(15 downto 0);
signal n21 : unsigned(15 downto 0);
signal n22 : unsigned(15 downto 0);
signal n23 : unsigned(15 downto 0);
signal n24 : unsigned(15 downto 0);
signal s25_1 : unsigned(15 downto 0);
signal s25_2 : unsigned(15 downto 0);
signal s26_1 : unsigned(0 downto 0);
signal s27_1 : unsigned(31 downto 0);
signal s28_1 : unsigned(0 downto 0);
signal s28_2 : unsigned(0 downto 0);
signal s28_3 : unsigned(31 downto 0);
signal s29_1 : unsigned(9 downto 0);
signal s29_2 : unsigned(0 downto 0);
component cf_fft_2048_8_7 is
port (
clock_c : in std_logic;
i1 : in  unsigned(15 downto 0);
i2 : in  unsigned(15 downto 0);
i3 : in  unsigned(0 downto 0);
i4 : in  unsigned(0 downto 0);
i5 : in  unsigned(0 downto 0);
o1 : out unsigned(15 downto 0);
o2 : out unsigned(15 downto 0));
end component cf_fft_2048_8_7;
component cf_fft_2048_8_35 is
port (
clock_c : in std_logic;
i1 : in  unsigned(1 downto 0);
i2 : in  unsigned(0 downto 0);
i3 : in  unsigned(0 downto 0);
o1 : out unsigned(0 downto 0));
end component cf_fft_2048_8_35;
component cf_fft_2048_8_31 is
port (
clock_c : in std_logic;
i1 : in  unsigned(31 downto 0);
i2 : in  unsigned(0 downto 0);
i3 : in  unsigned(8 downto 0);
i4 : in  unsigned(0 downto 0);
i5 : in  unsigned(0 downto 0);
i6 : in  unsigned(0 downto 0);
o1 : out unsigned(31 downto 0));
end component cf_fft_2048_8_31;
component cf_fft_2048_8_30 is
port (
clock_c : in std_logic;
i1 : in  unsigned(31 downto 0);
i2 : in  unsigned(0 downto 0);
i3 : in  unsigned(8 downto 0);
i4 : in  unsigned(0 downto 0);
i5 : in  unsigned(0 downto 0);
i6 : in  unsigned(0 downto 0);
o1 : out unsigned(0 downto 0);
o2 : out unsigned(0 downto 0);
o3 : out unsigned(31 downto 0));
end component cf_fft_2048_8_30;
component cf_fft_2048_8_26 is
port (
clock_c : in std_logic;
i1 : in  unsigned(0 downto 0);
i2 : in  unsigned(0 downto 0);
i3 : in  unsigned(0 downto 0);
o1 : out unsigned(9 downto 0);
o2 : out unsigned(0 downto 0));
end component cf_fft_2048_8_26;
begin
n1 <= s29_1(9 downto 9);
n2 <= s25_1 & s25_2;
process (clock_c) begin
  if rising_edge(clock_c) then
    if i5 = "1" then
      n3 <= "0";
    elsif i4 = "1" then
      n3 <= s29_2;
    end if;
  end if;
end process;
process (clock_c) begin
  if rising_edge(clock_c) then
    if i5 = "1" then
      n4 <= "0";
    elsif i4 = "1" then
      n4 <= n3;
    end if;
  end if;
end process;
process (clock_c) begin
  if rising_edge(clock_c) then
    if i5 = "1" then
      n5 <= "0";
    elsif i4 = "1" then
      n5 <= n4;
    end if;
  end if;
end process;
process (clock_c) begin
  if rising_edge(clock_c) then
    if i5 = "1" then
      n6 <= "0";
    elsif i4 = "1" then
      n6 <= n5;
    end if;
  end if;
end process;
n7 <= s29_1(9 downto 9) &
  s29_1(8 downto 8) &
  s29_1(7 downto 7) &
  s29_1(6 downto 6) &
  s29_1(5 downto 5) &
  s29_1(4 downto 4) &
  s29_1(3 downto 3) &
  s29_1(2 downto 2) &
  s29_1(1 downto 1);
process (clock_c) begin
  if rising_edge(clock_c) then
    if i5 = "1" then
      n8 <= "000000000";
    elsif i4 = "1" then
      n8 <= n7;
    end if;
  end if;
end process;
process (clock_c) begin
  if rising_edge(clock_c) then
    if i5 = "1" then
      n9 <= "000000000";
    elsif i4 = "1" then
      n9 <= n8;
    end if;
  end if;
end process;
process (clock_c) begin
  if rising_edge(clock_c) then
    if i5 = "1" then
      n10 <= "000000000";
    elsif i4 = "1" then
      n10 <= n9;
    end if;
  end if;
end process;
process (clock_c) begin
  if rising_edge(clock_c) then
    if i5 = "1" then
      n11 <= "000000000";
    elsif i4 = "1" then
      n11 <= n10;
    end if;
  end if;
end process;
n12 <= s29_1(0 downto 0);
process (clock_c) begin
  if rising_edge(clock_c) then
    if i5 = "1" then
      n13 <= "0";
    elsif i4 = "1" then
      n13 <= n12;
    end if;
  end if;
end process;
process (clock_c) begin
  if rising_edge(clock_c) then
    if i5 = "1" then
      n14 <= "0";
    elsif i4 = "1" then
      n14 <= n13;
    end if;
  end if;
end process;
process (clock_c) begin
  if rising_edge(clock_c) then
    if i5 = "1" then
      n15 <= "0";
    elsif i4 = "1" then
      n15 <= n14;
    end if;
  end if;
end process;
process (clock_c) begin
  if rising_edge(clock_c) then
    if i5 = "1" then
      n16 <= "0";
    elsif i4 = "1" then
      n16 <= n15;
    end if;
  end if;
end process;
n17 <= not n16;
n18 <= s28_2 & s28_1;
n19 <= s28_3(31 downto 31) &
  s28_3(30 downto 30) &
  s28_3(29 downto 29) &
  s28_3(28 downto 28) &
  s28_3(27 downto 27) &
  s28_3(26 downto 26) &
  s28_3(25 downto 25) &
  s28_3(24 downto 24) &
  s28_3(23 downto 23) &
  s28_3(22 downto 22) &
  s28_3(21 downto 21) &
  s28_3(20 downto 20) &
  s28_3(19 downto 19) &
  s28_3(18 downto 18) &
  s28_3(17 downto 17) &
  s28_3(16 downto 16);
n20 <= s28_3(15 downto 15) &
  s28_3(14 downto 14) &
  s28_3(13 downto 13) &
  s28_3(12 downto 12) &
  s28_3(11 downto 11) &
  s28_3(10 downto 10) &
  s28_3(9 downto 9) &
  s28_3(8 downto 8) &
  s28_3(7 downto 7) &
  s28_3(6 downto 6) &
  s28_3(5 downto 5) &
  s28_3(4 downto 4) &
  s28_3(3 downto 3) &
  s28_3(2 downto 2) &
  s28_3(1 downto 1) &
  s28_3(0 downto 0);
n21 <= s27_1(31 downto 31) &
  s27_1(30 downto 30) &
  s27_1(29 downto 29) &
  s27_1(28 downto 28) &
  s27_1(27 downto 27) &
  s27_1(26 downto 26) &
  s27_1(25 downto 25) &
  s27_1(24 downto 24) &
  s27_1(23 downto 23) &
  s27_1(22 downto 22) &
  s27_1(21 downto 21) &
  s27_1(20 downto 20) &
  s27_1(19 downto 19) &
  s27_1(18 downto 18) &
  s27_1(17 downto 17) &
  s27_1(16 downto 16);
n22 <= s27_1(15 downto 15) &
  s27_1(14 downto 14) &
  s27_1(13 downto 13) &
  s27_1(12 downto 12) &
  s27_1(11 downto 11) &
  s27_1(10 downto 10) &
  s27_1(9 downto 9) &
  s27_1(8 downto 8) &
  s27_1(7 downto 7) &
  s27_1(6 downto 6) &
  s27_1(5 downto 5) &
  s27_1(4 downto 4) &
  s27_1(3 downto 3) &
  s27_1(2 downto 2) &
  s27_1(1 downto 1) &
  s27_1(0 downto 0);
n23 <= n20 when s26_1 = "1" else n19;
n24 <= n22 when s26_1 = "1" else n21;
s25 : cf_fft_2048_8_7 port map (clock_c, i2, i3, n1, i4, i5, s25_1, s25_2);
s26 : cf_fft_2048_8_35 port map (clock_c, n18, i4, i5, s26_1);
s27 : cf_fft_2048_8_31 port map (clock_c, n2, n6, n11, n16, i4, i5, s27_1);
s28 : cf_fft_2048_8_30 port map (clock_c, n2, n6, n11, n17, i4, i5, s28_1, s28_2, s28_3);
s29 : cf_fft_2048_8_26 port map (clock_c, i1, i4, i5, s29_1, s29_2);
o3 <= n24;
o2 <= n23;
o1 <= s28_1;
end architecture rtl;

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
entity cf_fft_2048_8_5 is
port (
clock_c : in std_logic;
i1 : in  unsigned(0 downto 0);
i2 : in  unsigned(15 downto 0);
i3 : in  unsigned(15 downto 0);
i4 : in  unsigned(0 downto 0);
i5 : in  unsigned(0 downto 0);
o1 : out unsigned(0 downto 0);
o2 : out unsigned(15 downto 0);
o3 : out unsigned(15 downto 0));
end entity cf_fft_2048_8_5;
architecture rtl of cf_fft_2048_8_5 is
signal n1 : unsigned(0 downto 0);
signal n2 : unsigned(31 downto 0);
signal n3 : unsigned(0 downto 0) := "0";
signal n4 : unsigned(0 downto 0) := "0";
signal n5 : unsigned(0 downto 0) := "0";
signal n6 : unsigned(0 downto 0) := "0";
signal n7 : unsigned(8 downto 0);
signal n8 : unsigned(8 downto 0) := "000000000";
signal n9 : unsigned(8 downto 0) := "000000000";
signal n10 : unsigned(8 downto 0) := "000000000";
signal n11 : unsigned(8 downto 0) := "000000000";
signal n12 : unsigned(0 downto 0);
signal n13 : unsigned(0 downto 0) := "0";
signal n14 : unsigned(0 downto 0) := "0";
signal n15 : unsigned(0 downto 0) := "0";
signal n16 : unsigned(0 downto 0) := "0";
signal n17 : unsigned(0 downto 0);
signal n18 : unsigned(1 downto 0);
signal n19 : unsigned(15 downto 0);
signal n20 : unsigned(15 downto 0);
signal n21 : unsigned(15 downto 0);
signal n22 : unsigned(15 downto 0);
signal n23 : unsigned(15 downto 0);
signal n24 : unsigned(15 downto 0);
signal s25_1 : unsigned(15 downto 0);
signal s25_2 : unsigned(15 downto 0);
signal s26_1 : unsigned(0 downto 0);
signal s27_1 : unsigned(31 downto 0);
signal s28_1 : unsigned(0 downto 0);
signal s28_2 : unsigned(0 downto 0);
signal s28_3 : unsigned(31 downto 0);
signal s29_1 : unsigned(9 downto 0);
signal s29_2 : unsigned(0 downto 0);
component cf_fft_2048_8_7 is
port (
clock_c : in std_logic;
i1 : in  unsigned(15 downto 0);
i2 : in  unsigned(15 downto 0);
i3 : in  unsigned(0 downto 0);
i4 : in  unsigned(0 downto 0);
i5 : in  unsigned(0 downto 0);
o1 : out unsigned(15 downto 0);
o2 : out unsigned(15 downto 0));
end component cf_fft_2048_8_7;
component cf_fft_2048_8_35 is
port (
clock_c : in std_logic;
i1 : in  unsigned(1 downto 0);
i2 : in  unsigned(0 downto 0);
i3 : in  unsigned(0 downto 0);
o1 : out unsigned(0 downto 0));
end component cf_fft_2048_8_35;
component cf_fft_2048_8_31 is
port (
clock_c : in std_logic;
i1 : in  unsigned(31 downto 0);
i2 : in  unsigned(0 downto 0);
i3 : in  unsigned(8 downto 0);
i4 : in  unsigned(0 downto 0);
i5 : in  unsigned(0 downto 0);
i6 : in  unsigned(0 downto 0);
o1 : out unsigned(31 downto 0));
end component cf_fft_2048_8_31;
component cf_fft_2048_8_30 is
port (
clock_c : in std_logic;
i1 : in  unsigned(31 downto 0);
i2 : in  unsigned(0 downto 0);
i3 : in  unsigned(8 downto 0);
i4 : in  unsigned(0 downto 0);
i5 : in  unsigned(0 downto 0);
i6 : in  unsigned(0 downto 0);
o1 : out unsigned(0 downto 0);
o2 : out unsigned(0 downto 0);
o3 : out unsigned(31 downto 0));
end component cf_fft_2048_8_30;
component cf_fft_2048_8_26 is
port (
clock_c : in std_logic;
i1 : in  unsigned(0 downto 0);
i2 : in  unsigned(0 downto 0);
i3 : in  unsigned(0 downto 0);
o1 : out unsigned(9 downto 0);
o2 : out unsigned(0 downto 0));
end component cf_fft_2048_8_26;
begin
n1 <= "0";
n2 <= s25_1 & s25_2;
process (clock_c) begin
  if rising_edge(clock_c) then
    if i5 = "1" then
      n3 <= "0";
    elsif i4 = "1" then
      n3 <= s29_2;
    end if;
  end if;
end process;
process (clock_c) begin
  if rising_edge(clock_c) then
    if i5 = "1" then
      n4 <= "0";
    elsif i4 = "1" then
      n4 <= n3;
    end if;
  end if;
end process;
process (clock_c) begin
  if rising_edge(clock_c) then
    if i5 = "1" then
      n5 <= "0";
    elsif i4 = "1" then
      n5 <= n4;
    end if;
  end if;
end process;
process (clock_c) begin
  if rising_edge(clock_c) then
    if i5 = "1" then
      n6 <= "0";
    elsif i4 = "1" then
      n6 <= n5;
    end if;
  end if;
end process;
n7 <= s29_1(9 downto 9) &
  s29_1(8 downto 8) &
  s29_1(7 downto 7) &
  s29_1(6 downto 6) &
  s29_1(5 downto 5) &
  s29_1(4 downto 4) &
  s29_1(3 downto 3) &
  s29_1(2 downto 2) &
  s29_1(1 downto 1);
process (clock_c) begin
  if rising_edge(clock_c) then
    if i5 = "1" then
      n8 <= "000000000";
    elsif i4 = "1" then
      n8 <= n7;
    end if;
  end if;
end process;
process (clock_c) begin
  if rising_edge(clock_c) then
    if i5 = "1" then
      n9 <= "000000000";
    elsif i4 = "1" then
      n9 <= n8;
    end if;
  end if;
end process;
process (clock_c) begin
  if rising_edge(clock_c) then
    if i5 = "1" then
      n10 <= "000000000";
    elsif i4 = "1" then
      n10 <= n9;
    end if;
  end if;
end process;
process (clock_c) begin
  if rising_edge(clock_c) then
    if i5 = "1" then
      n11 <= "000000000";
    elsif i4 = "1" then
      n11 <= n10;
    end if;
  end if;
end process;
n12 <= s29_1(0 downto 0);
process (clock_c) begin
  if rising_edge(clock_c) then
    if i5 = "1" then
      n13 <= "0";
    elsif i4 = "1" then
      n13 <= n12;
    end if;
  end if;
end process;
process (clock_c) begin
  if rising_edge(clock_c) then
    if i5 = "1" then
      n14 <= "0";
    elsif i4 = "1" then
      n14 <= n13;
    end if;
  end if;
end process;
process (clock_c) begin
  if rising_edge(clock_c) then
    if i5 = "1" then
      n15 <= "0";
    elsif i4 = "1" then
      n15 <= n14;
    end if;
  end if;
end process;
process (clock_c) begin
  if rising_edge(clock_c) then
    if i5 = "1" then
      n16 <= "0";
    elsif i4 = "1" then
      n16 <= n15;
    end if;
  end if;
end process;
n17 <= not n16;
n18 <= s28_2 & s28_1;
n19 <= s28_3(31 downto 31) &
  s28_3(30 downto 30) &
  s28_3(29 downto 29) &
  s28_3(28 downto 28) &
  s28_3(27 downto 27) &
  s28_3(26 downto 26) &
  s28_3(25 downto 25) &
  s28_3(24 downto 24) &
  s28_3(23 downto 23) &
  s28_3(22 downto 22) &
  s28_3(21 downto 21) &
  s28_3(20 downto 20) &
  s28_3(19 downto 19) &
  s28_3(18 downto 18) &
  s28_3(17 downto 17) &
  s28_3(16 downto 16);
n20 <= s28_3(15 downto 15) &
  s28_3(14 downto 14) &
  s28_3(13 downto 13) &
  s28_3(12 downto 12) &
  s28_3(11 downto 11) &
  s28_3(10 downto 10) &
  s28_3(9 downto 9) &
  s28_3(8 downto 8) &
  s28_3(7 downto 7) &
  s28_3(6 downto 6) &
  s28_3(5 downto 5) &
  s28_3(4 downto 4) &
  s28_3(3 downto 3) &
  s28_3(2 downto 2) &
  s28_3(1 downto 1) &
  s28_3(0 downto 0);
n21 <= s27_1(31 downto 31) &
  s27_1(30 downto 30) &
  s27_1(29 downto 29) &
  s27_1(28 downto 28) &
  s27_1(27 downto 27) &
  s27_1(26 downto 26) &
  s27_1(25 downto 25) &
  s27_1(24 downto 24) &
  s27_1(23 downto 23) &
  s27_1(22 downto 22) &
  s27_1(21 downto 21) &
  s27_1(20 downto 20) &
  s27_1(19 downto 19) &
  s27_1(18 downto 18) &
  s27_1(17 downto 17) &
  s27_1(16 downto 16);
n22 <= s27_1(15 downto 15) &
  s27_1(14 downto 14) &
  s27_1(13 downto 13) &
  s27_1(12 downto 12) &
  s27_1(11 downto 11) &
  s27_1(10 downto 10) &
  s27_1(9 downto 9) &
  s27_1(8 downto 8) &
  s27_1(7 downto 7) &
  s27_1(6 downto 6) &
  s27_1(5 downto 5) &
  s27_1(4 downto 4) &
  s27_1(3 downto 3) &
  s27_1(2 downto 2) &
  s27_1(1 downto 1) &
  s27_1(0 downto 0);
n23 <= n20 when s26_1 = "1" else n19;
n24 <= n22 when s26_1 = "1" else n21;
s25 : cf_fft_2048_8_7 port map (clock_c, i2, i3, n1, i4, i5, s25_1, s25_2);
s26 : cf_fft_2048_8_35 port map (clock_c, n18, i4, i5, s26_1);
s27 : cf_fft_2048_8_31 port map (clock_c, n2, n6, n11, n16, i4, i5, s27_1);
s28 : cf_fft_2048_8_30 port map (clock_c, n2, n6, n11, n17, i4, i5, s28_1, s28_2, s28_3);
s29 : cf_fft_2048_8_26 port map (clock_c, i1, i4, i5, s29_1, s29_2);
o3 <= n24;
o2 <= n23;
o1 <= s28_1;
end architecture rtl;

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
entity cf_fft_2048_8_4 is
port (
clock_c : in std_logic;
i1 : in  unsigned(0 downto 0);
i2 : in  unsigned(31 downto 0);
i3 : in  unsigned(0 downto 0);
i4 : in  unsigned(8 downto 0);
i5 : in  unsigned(0 downto 0);
i6 : in  unsigned(0 downto 0);
o1 : out unsigned(31 downto 0));
end entity cf_fft_2048_8_4;
architecture rtl of cf_fft_2048_8_4 is
signal n1 : unsigned(8 downto 0);
signal n2 : unsigned(8 downto 0);
signal n3 : unsigned(8 downto 0) := "000000000";
signal n4 : unsigned(0 downto 0);
signal n5 : unsigned(0 downto 0);
signal n6 : unsigned(31 downto 0);
signal n6a : unsigned(8 downto 0) := "000000000";
type   n6mt is array (511 downto 0) of unsigned(31 downto 0);
signal n6m : n6mt;
signal n7 : unsigned(0 downto 0);
signal n8 : unsigned(31 downto 0);
signal n8a : unsigned(8 downto 0) := "000000000";
type   n8mt is array (511 downto 0) of unsigned(31 downto 0);
signal n8m : n8mt;
signal n9 : unsigned(0 downto 0) := "0";
signal n10 : unsigned(31 downto 0);
signal n11 : unsigned(0 downto 0);
signal s12_1 : unsigned(0 downto 0);
component cf_fft_2048_8_32 is
port (
clock_c : in std_logic;
i1 : in  unsigned(0 downto 0);
i2 : in  unsigned(0 downto 0);
i3 : in  unsigned(0 downto 0);
o1 : out unsigned(0 downto 0));
end component cf_fft_2048_8_32;
begin
n1 <= "000000001";
n2 <= n3 + n1;
process (clock_c) begin
  if rising_edge(clock_c) then
    if n11 = "1" then
      n3 <= "000000000";
    elsif i5 = "1" then
      n3 <= n2;
    end if;
  end if;
end process;
n4 <= not s12_1;
n5 <= i3 and n4;
process (clock_c) begin
  if rising_edge(clock_c) then
    if i5 = "1" then
      if n5 = "1" then
        n6m(to_integer(i4)) <= i2;
      end if;
      n6a <= n3;
    end if;
  end if;
end process;
n6 <= n6m(to_integer(n6a));
n7 <= i3 and s12_1;
process (clock_c) begin
  if rising_edge(clock_c) then
    if i5 = "1" then
      if n7 = "1" then
        n8m(to_integer(i4)) <= i2;
      end if;
      n8a <= n3;
    end if;
  end if;
end process;
n8 <= n8m(to_integer(n8a));
process (clock_c) begin
  if rising_edge(clock_c) then
    if i6 = "1" then
      n9 <= "0";
    elsif i5 = "1" then
      n9 <= n4;
    end if;
  end if;
end process;
n10 <= n8 when n9 = "1" else n6;
n11 <= i1 or i6;
s12 : cf_fft_2048_8_32 port map (clock_c, i1, i5, i6, s12_1);
o1 <= n10;
end architecture rtl;

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
entity cf_fft_2048_8_3 is
port (
clock_c : in std_logic;
i1 : in  unsigned(0 downto 0);
i2 : in  unsigned(31 downto 0);
i3 : in  unsigned(0 downto 0);
i4 : in  unsigned(8 downto 0);
i5 : in  unsigned(0 downto 0);
i6 : in  unsigned(0 downto 0);
o1 : out unsigned(0 downto 0);
o2 : out unsigned(0 downto 0);
o3 : out unsigned(31 downto 0));
end entity cf_fft_2048_8_3;
architecture rtl of cf_fft_2048_8_3 is
signal n1 : unsigned(8 downto 0);
signal n2 : unsigned(8 downto 0);
signal n3 : unsigned(8 downto 0) := "000000000";
signal n4 : unsigned(0 downto 0);
signal n5 : unsigned(0 downto 0) := "0";
signal n6 : unsigned(8 downto 0);
signal n7 : unsigned(0 downto 0);
signal n8 : unsigned(0 downto 0);
signal n9 : unsigned(31 downto 0);
signal n9a : unsigned(8 downto 0) := "000000000";
type   n9mt is array (511 downto 0) of unsigned(31 downto 0);
signal n9m : n9mt;
signal n10 : unsigned(0 downto 0);
signal n11 : unsigned(31 downto 0);
signal n11a : unsigned(8 downto 0) := "000000000";
type   n11mt is array (511 downto 0) of unsigned(31 downto 0);
signal n11m : n11mt;
signal n12 : unsigned(0 downto 0) := "0";
signal n13 : unsigned(31 downto 0);
signal n14 : unsigned(0 downto 0);
signal s15_1 : unsigned(0 downto 0);
component cf_fft_2048_8_32 is
port (
clock_c : in std_logic;
i1 : in  unsigned(0 downto 0);
i2 : in  unsigned(0 downto 0);
i3 : in  unsigned(0 downto 0);
o1 : out unsigned(0 downto 0));
end component cf_fft_2048_8_32;
begin
n1 <= "000000001";
n2 <= n3 + n1;
process (clock_c) begin
  if rising_edge(clock_c) then
    if n14 = "1" then
      n3 <= "000000000";
    elsif i5 = "1" then
      n3 <= n2;
    end if;
  end if;
end process;
n4 <= not s15_1;
process (clock_c) begin
  if rising_edge(clock_c) then
    if i6 = "1" then
      n5 <= "0";
    elsif i5 = "1" then
      n5 <= i1;
    end if;
  end if;
end process;
n6 <= "000000000";
n7 <= "1" when n3 = n6 else "0";
n8 <= i3 and n4;
process (clock_c) begin
  if rising_edge(clock_c) then
    if i5 = "1" then
      if n8 = "1" then
        n9m(to_integer(i4)) <= i2;
      end if;
      n9a <= n3;
    end if;
  end if;
end process;
n9 <= n9m(to_integer(n9a));
n10 <= i3 and s15_1;
process (clock_c) begin
  if rising_edge(clock_c) then
    if i5 = "1" then
      if n10 = "1" then
        n11m(to_integer(i4)) <= i2;
      end if;
      n11a <= n3;
    end if;
  end if;
end process;
n11 <= n11m(to_integer(n11a));
process (clock_c) begin
  if rising_edge(clock_c) then
    if i6 = "1" then
      n12 <= "0";
    elsif i5 = "1" then
      n12 <= n4;
    end if;
  end if;
end process;
n13 <= n11 when n12 = "1" else n9;
n14 <= i1 or i6;
s15 : cf_fft_2048_8_32 port map (clock_c, i1, i5, i6, s15_1);
o3 <= n13;
o2 <= n7;
o1 <= n5;
end architecture rtl;

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
entity cf_fft_2048_8_2 is
port (
clock_c : in std_logic;
i1 : in  unsigned(0 downto 0);
i2 : in  unsigned(15 downto 0);
i3 : in  unsigned(15 downto 0);
i4 : in  unsigned(0 downto 0);
i5 : in  unsigned(0 downto 0);
o1 : out unsigned(0 downto 0);
o2 : out unsigned(15 downto 0);
o3 : out unsigned(15 downto 0));
end entity cf_fft_2048_8_2;
architecture rtl of cf_fft_2048_8_2 is
signal n1 : unsigned(31 downto 0);
signal n2 : unsigned(0 downto 0);
signal n3 : unsigned(0 downto 0);
signal n4 : unsigned(8 downto 0);
signal n5 : unsigned(8 downto 0);
signal n6 : unsigned(1 downto 0);
signal n7 : unsigned(15 downto 0);
signal n8 : unsigned(15 downto 0);
signal n9 : unsigned(15 downto 0);
signal n10 : unsigned(15 downto 0);
signal n11 : unsigned(15 downto 0);
signal n12 : unsigned(15 downto 0);
signal s13_1 : unsigned(0 downto 0);
signal s14_1 : unsigned(31 downto 0);
signal s15_1 : unsigned(0 downto 0);
signal s15_2 : unsigned(0 downto 0);
signal s15_3 : unsigned(31 downto 0);
signal s16_1 : unsigned(9 downto 0);
signal s16_2 : unsigned(0 downto 0);
component cf_fft_2048_8_35 is
port (
clock_c : in std_logic;
i1 : in  unsigned(1 downto 0);
i2 : in  unsigned(0 downto 0);
i3 : in  unsigned(0 downto 0);
o1 : out unsigned(0 downto 0));
end component cf_fft_2048_8_35;
component cf_fft_2048_8_4 is
port (
clock_c : in std_logic;
i1 : in  unsigned(0 downto 0);
i2 : in  unsigned(31 downto 0);
i3 : in  unsigned(0 downto 0);
i4 : in  unsigned(8 downto 0);
i5 : in  unsigned(0 downto 0);
i6 : in  unsigned(0 downto 0);
o1 : out unsigned(31 downto 0));
end component cf_fft_2048_8_4;
component cf_fft_2048_8_3 is
port (
clock_c : in std_logic;
i1 : in  unsigned(0 downto 0);
i2 : in  unsigned(31 downto 0);
i3 : in  unsigned(0 downto 0);
i4 : in  unsigned(8 downto 0);
i5 : in  unsigned(0 downto 0);
i6 : in  unsigned(0 downto 0);
o1 : out unsigned(0 downto 0);
o2 : out unsigned(0 downto 0);
o3 : out unsigned(31 downto 0));
end component cf_fft_2048_8_3;
component cf_fft_2048_8_26 is
port (
clock_c : in std_logic;
i1 : in  unsigned(0 downto 0);
i2 : in  unsigned(0 downto 0);
i3 : in  unsigned(0 downto 0);
o1 : out unsigned(9 downto 0);
o2 : out unsigned(0 downto 0));
end component cf_fft_2048_8_26;
begin
n1 <= i2 & i3;
n2 <= s16_1(9 downto 9);
n3 <= not n2;
n4 <= s16_1(8 downto 8) &
  s16_1(7 downto 7) &
  s16_1(6 downto 6) &
  s16_1(5 downto 5) &
  s16_1(4 downto 4) &
  s16_1(3 downto 3) &
  s16_1(2 downto 2) &
  s16_1(1 downto 1) &
  s16_1(0 downto 0);
n5 <= n4(0 downto 0) &
  n4(1 downto 1) &
  n4(2 downto 2) &
  n4(3 downto 3) &
  n4(4 downto 4) &
  n4(5 downto 5) &
  n4(6 downto 6) &
  n4(7 downto 7) &
  n4(8 downto 8);
n6 <= s15_2 & s15_1;
n7 <= s15_3(31 downto 31) &
  s15_3(30 downto 30) &
  s15_3(29 downto 29) &
  s15_3(28 downto 28) &
  s15_3(27 downto 27) &
  s15_3(26 downto 26) &
  s15_3(25 downto 25) &
  s15_3(24 downto 24) &
  s15_3(23 downto 23) &
  s15_3(22 downto 22) &
  s15_3(21 downto 21) &
  s15_3(20 downto 20) &
  s15_3(19 downto 19) &
  s15_3(18 downto 18) &
  s15_3(17 downto 17) &
  s15_3(16 downto 16);
n8 <= s15_3(15 downto 15) &
  s15_3(14 downto 14) &
  s15_3(13 downto 13) &
  s15_3(12 downto 12) &
  s15_3(11 downto 11) &
  s15_3(10 downto 10) &
  s15_3(9 downto 9) &
  s15_3(8 downto 8) &
  s15_3(7 downto 7) &
  s15_3(6 downto 6) &
  s15_3(5 downto 5) &
  s15_3(4 downto 4) &
  s15_3(3 downto 3) &
  s15_3(2 downto 2) &
  s15_3(1 downto 1) &
  s15_3(0 downto 0);
n9 <= s14_1(31 downto 31) &
  s14_1(30 downto 30) &
  s14_1(29 downto 29) &
  s14_1(28 downto 28) &
  s14_1(27 downto 27) &
  s14_1(26 downto 26) &
  s14_1(25 downto 25) &
  s14_1(24 downto 24) &
  s14_1(23 downto 23) &
  s14_1(22 downto 22) &
  s14_1(21 downto 21) &
  s14_1(20 downto 20) &
  s14_1(19 downto 19) &
  s14_1(18 downto 18) &
  s14_1(17 downto 17) &
  s14_1(16 downto 16);
n10 <= s14_1(15 downto 15) &
  s14_1(14 downto 14) &
  s14_1(13 downto 13) &
  s14_1(12 downto 12) &
  s14_1(11 downto 11) &
  s14_1(10 downto 10) &
  s14_1(9 downto 9) &
  s14_1(8 downto 8) &
  s14_1(7 downto 7) &
  s14_1(6 downto 6) &
  s14_1(5 downto 5) &
  s14_1(4 downto 4) &
  s14_1(3 downto 3) &
  s14_1(2 downto 2) &
  s14_1(1 downto 1) &
  s14_1(0 downto 0);
n11 <= n8 when s13_1 = "1" else n7;
n12 <= n10 when s13_1 = "1" else n9;
s13 : cf_fft_2048_8_35 port map (clock_c, n6, i4, i5, s13_1);
s14 : cf_fft_2048_8_4 port map (clock_c, s16_2, n1, n2, n5, i4, i5, s14_1);
s15 : cf_fft_2048_8_3 port map (clock_c, s16_2, n1, n3, n5, i4, i5, s15_1, s15_2, s15_3);
s16 : cf_fft_2048_8_26 port map (clock_c, i1, i4, i5, s16_1, s16_2);
o3 <= n12;
o2 <= n11;
o1 <= s15_1;
end architecture rtl;

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
entity cf_fft_2048_8_1 is
port (
clock_c : in std_logic;
i1 : in  unsigned(0 downto 0);
i2 : in  unsigned(15 downto 0);
i3 : in  unsigned(15 downto 0);
i4 : in  unsigned(0 downto 0);
i5 : in  unsigned(0 downto 0);
o1 : out unsigned(0 downto 0);
o2 : out unsigned(15 downto 0);
o3 : out unsigned(15 downto 0));
end entity cf_fft_2048_8_1;
architecture rtl of cf_fft_2048_8_1 is
signal s1_1 : unsigned(0 downto 0);
signal s1_2 : unsigned(15 downto 0);
signal s1_3 : unsigned(15 downto 0);
signal s2_1 : unsigned(0 downto 0);
signal s2_2 : unsigned(15 downto 0);
signal s2_3 : unsigned(15 downto 0);
signal s3_1 : unsigned(0 downto 0);
signal s3_2 : unsigned(15 downto 0);
signal s3_3 : unsigned(15 downto 0);
signal s4_1 : unsigned(0 downto 0);
signal s4_2 : unsigned(15 downto 0);
signal s4_3 : unsigned(15 downto 0);
signal s5_1 : unsigned(0 downto 0);
signal s5_2 : unsigned(15 downto 0);
signal s5_3 : unsigned(15 downto 0);
component cf_fft_2048_8_25 is
port (
clock_c : in std_logic;
i1 : in  unsigned(0 downto 0);
i2 : in  unsigned(15 downto 0);
i3 : in  unsigned(15 downto 0);
i4 : in  unsigned(0 downto 0);
i5 : in  unsigned(0 downto 0);
o1 : out unsigned(0 downto 0);
o2 : out unsigned(15 downto 0);
o3 : out unsigned(15 downto 0));
end component cf_fft_2048_8_25;
component cf_fft_2048_8_8 is
port (
clock_c : in std_logic;
i1 : in  unsigned(0 downto 0);
i2 : in  unsigned(15 downto 0);
i3 : in  unsigned(15 downto 0);
i4 : in  unsigned(0 downto 0);
i5 : in  unsigned(0 downto 0);
o1 : out unsigned(0 downto 0);
o2 : out unsigned(15 downto 0);
o3 : out unsigned(15 downto 0));
end component cf_fft_2048_8_8;
component cf_fft_2048_8_6 is
port (
clock_c : in std_logic;
i1 : in  unsigned(0 downto 0);
i2 : in  unsigned(15 downto 0);
i3 : in  unsigned(15 downto 0);
i4 : in  unsigned(0 downto 0);
i5 : in  unsigned(0 downto 0);
o1 : out unsigned(0 downto 0);
o2 : out unsigned(15 downto 0);
o3 : out unsigned(15 downto 0));
end component cf_fft_2048_8_6;
component cf_fft_2048_8_5 is
port (
clock_c : in std_logic;
i1 : in  unsigned(0 downto 0);
i2 : in  unsigned(15 downto 0);
i3 : in  unsigned(15 downto 0);
i4 : in  unsigned(0 downto 0);
i5 : in  unsigned(0 downto 0);
o1 : out unsigned(0 downto 0);
o2 : out unsigned(15 downto 0);
o3 : out unsigned(15 downto 0));
end component cf_fft_2048_8_5;
component cf_fft_2048_8_2 is
port (
clock_c : in std_logic;
i1 : in  unsigned(0 downto 0);
i2 : in  unsigned(15 downto 0);
i3 : in  unsigned(15 downto 0);
i4 : in  unsigned(0 downto 0);
i5 : in  unsigned(0 downto 0);
o1 : out unsigned(0 downto 0);
o2 : out unsigned(15 downto 0);
o3 : out unsigned(15 downto 0));
end component cf_fft_2048_8_2;
begin
s1 : cf_fft_2048_8_25 port map (clock_c, s3_1, s3_2, s3_3, i4, i5, s1_1, s1_2, s1_3);
s2 : cf_fft_2048_8_8 port map (clock_c, s1_1, s1_2, s1_3, i4, i5, s2_1, s2_2, s2_3);
s3 : cf_fft_2048_8_6 port map (clock_c, s4_1, s4_2, s4_3, i4, i5, s3_1, s3_2, s3_3);
s4 : cf_fft_2048_8_5 port map (clock_c, s5_1, s5_2, s5_3, i4, i5, s4_1, s4_2, s4_3);
s5 : cf_fft_2048_8_2 port map (clock_c, i1, i2, i3, i4, i5, s5_1, s5_2, s5_3);
o3 <= s2_3;
o2 <= s2_2;
o1 <= s2_1;
end architecture rtl;

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
entity cf_fft_2048_8 is
port(
signal clock_c : in std_logic;
signal enable_i : in unsigned(0 downto 0);
signal reset_i : in unsigned(0 downto 0);
signal sync_i : in unsigned(0 downto 0);
signal data_0_i : in unsigned(15 downto 0);
signal data_1_i : in unsigned(15 downto 0);
signal sync_o : out unsigned(0 downto 0);
signal data_0_o : out unsigned(15 downto 0);
signal data_1_o : out unsigned(15 downto 0));
end entity cf_fft_2048_8;
architecture rtl of cf_fft_2048_8 is
component cf_fft_2048_8_1 is
port (
clock_c : in std_logic;
i1 : in  unsigned(0 downto 0);
i2 : in  unsigned(15 downto 0);
i3 : in  unsigned(15 downto 0);
i4 : in  unsigned(0 downto 0);
i5 : in  unsigned(0 downto 0);
o1 : out unsigned(0 downto 0);
o2 : out unsigned(15 downto 0);
o3 : out unsigned(15 downto 0));
end component cf_fft_2048_8_1;
signal n1 : unsigned(0 downto 0);
signal n2 : unsigned(15 downto 0);
signal n3 : unsigned(15 downto 0);
begin
s1 : cf_fft_2048_8_1 port map (clock_c, sync_i, data_0_i, data_1_i, enable_i, reset_i, n1, n2, n3);
sync_o <= n1;
data_0_o <= n2;
data_1_o <= n3;
end architecture rtl;


